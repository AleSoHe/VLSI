* FLIP FLOP LAYOUT LEVEL

.options POST=1 parhier=local

.subckt flip-flop c cn d q rn
cg3303 532:vdd gnd  c=4.80879e-16
c3302 532:vdd x12|src  c=1.11383e-19
c3301 532:vdd 259:4  c=1.46892e-17
c3300 532:vdd 303:2  c=1.17625e-18
c3299 532:vdd 246:4  c=1.03155e-17
c3298 532:vdd 433:3  c=2.50243e-18
c3297 532:vdd 426:3  c=1.50108e-17
c3296 532:vdd 147:16  c=4.79229e-17
c3295 532:vdd 427:3  c=3.13789e-18
c3294 532:vdd 151:16  c=4.85048e-17
c3293 532:vdd 425:3  c=1.59881e-17
c3292 532:vdd x17|drn  c=2.81188e-20
c3291 532:vdd 218:9  c=2.59473e-18
c3290 532:vdd 305:2  c=1.53055e-18
c3289 532:vdd 306:2  c=2.13918e-17
c3288 532:vdd 350:2  c=1.71922e-17
c3287 532:vdd 319:2  c=1.49018e-17
c3286 532:vdd 307:2  c=9.95111e-18
c3285 532:vdd 135:14  c=4.43255e-17
c3284 532:vdd 65:d  c=1.15209e-18
c3283 532:vdd 61:d  c=1.58855e-18
c3282 532:vdd 32:rn  c=1.21259e-17
c3281 532:vdd 220:9  c=2.81847e-18
c3280 532:vdd x21|src  c=7.18097e-20
c3279 532:vdd 71:d  c=1.15209e-18
c3278 532:vdd 56:d  c=1.17806e-18
c3277 532:vdd x24|drn  c=1.25725e-19
c3276 532:vdd x24|src  c=7.43815e-20
c3275 532:vdd x25|drn  c=1.32484e-19
c3274 532:vdd 58:d  c=1.95271e-19
c3273 532:vdd x26|src  c=1.21582e-19
c3272 532:vdd 138:14  c=3.43404e-18
c3271 532:vdd x28|drn  c=1.03775e-19
c3270 532:vdd 329:2  c=3.27894e-18
c3269 532:vdd 140:14  c=3.44336e-18
c3268 532:vdd 167:16  c=2.53283e-18
c3267 532:vdd 281:4  c=4.15716e-19
c3266 532:vdd 157:16  c=4.03017e-17
c3265 532:vdd 266:4  c=1.83324e-18
c3264 532:vdd 292:4  c=1.15216e-18
c3263 532:vdd 143:14  c=2.94844e-18
c3262 532:vdd 48:rn  c=9.412e-19
c3261 532:vdd 289:4  c=5.27991e-17
c3260 532:vdd 202:9  c=4.34005e-17
c3259 532:vdd 169:16  c=2.60107e-18
c3258 532:vdd 33:rn  c=1.92844e-18
c3257 532:vdd 293:4  c=5.16879e-17
c3256 532:vdd 239:9  c=4.49308e-17
c3255 532:vdd 23:rn  c=1.92844e-18
c3254 532:vdd 247:4  c=2.59023e-19
c3253 532:vdd 420:cn  c=1.20758e-20
c3252 532:vdd 338:2  c=4.90469e-17
c3251 532:vdd 310:2  c=3.86408e-18
c3250 532:vdd 171:16  c=3.45659e-18
c3249 532:vdd 434:3  c=5.4153e-17
c3248 532:vdd gnd  c=7.32059e-21
c3247 532:vdd 49:rn  c=1.92844e-18
c3246 532:vdd 51:rn  c=1.70517e-19
c3245 532:vdd 237:9  c=1.03551e-18
c3244 532:vdd 4:rn  c=1.6265e-18
c3243 532:vdd 435:3  c=5.55286e-17
c3242 532:vdd 354:cn  c=1.70601e-18
c3241 532:vdd 240:9  c=4.7011e-17
c3240 532:vdd 206:9  c=6.19196e-18
c3239 532:vdd 337:2  c=4.29494e-20
c3238 532:vdd 412:cn  c=1.82034e-18
c3237 532:vdd 353:2  c=1.33975e-18
c3236 532:vdd 367:cn  c=8.99218e-19
c3235 532:vdd 311:2  c=1.48594e-18
c3234 532:vdd 390:cn  c=2.83115e-18
c3233 532:vdd 347:2  c=5.27286e-17
c3232 532:vdd 136:14  c=4.93046e-17
c3231 532:vdd 352:2  c=5.14341e-17
c3230 532:vdd m10|x1|gate  c=4.80249e-19
c3229 532:vdd 208:9  c=2.77182e-18
c3228 532:vdd m10|x1|src  c=8.67494e-20
c3227 532:vdd 198:9  c=4.69608e-17
c3226 532:vdd 392:cn  c=1.81037e-18
c3225 532:vdd 144:14  c=4.789e-17
c3224 532:vdd m11|x1|drn  c=9.33909e-20
c3223 532:vdd m11|x1|gate  c=6.08998e-19
c3222 532:vdd m11|x1|src  c=9.00999e-20
c3221 532:vdd m18|x1|bulk  c=2.71746e-16
c3220 532:vdd 269:4  c=2.60889e-18
c3219 532:vdd 242:4  c=1.09387e-18
c3218 532:vdd 252:4  c=2.39037e-18
c3217 532:vdd 40:rn  c=1.64677e-18
c3216 532:vdd 216:9  c=2.60107e-18
c3215 532:vdd 230:9  c=1.03701e-18
c3214 532:vdd 322:2  c=2.64455e-18
c3213 532:vdd 232:9  c=1.44432e-19
c3212 532:vdd 339:2  c=1.15091e-18
c3211 532:vdd x10|drn  c=9.48935e-20
c3210 532:vdd 50:rn  c=1.53286e-18
c3209 532:vdd 312:2  c=3.22513e-18
c3208 532:vdd 340:2  c=1.83143e-18
c3207 532:vdd 431:3  c=3.38322e-18
c3206 532:vdd 294:4  c=1.63412e-17
c3205 532:vdd 351:2  c=1.15091e-18
cg3204 x30|src gnd  c=1.76057e-20
c3203 x30|src 144:14  c=2.36627e-19
c3202 x30|src 71:d  c=7.43977e-19
c3201 x30|src 364:cn  c=4.19174e-20
c3200 x30|src 58:d  c=6.47761e-19
c3199 x30|src 143:14  c=7.76216e-19
c3198 x30|src 64:d  c=7.43977e-19
c3197 x30|src gnd  c=8.65274e-20
c3196 x29|src 437:gnd  c=7.09333e-20
c3195 x29|src 306:2  c=5.48108e-19
c3194 x29|src 351:2  c=6.97626e-19
c3193 x29|src 220:9  c=7.76216e-19
c3192 x29|src 328:2  c=6.97626e-19
c3191 x29|src 364:cn  c=1.01633e-20
c3190 x29|src 308:2  c=1.19594e-19
c3189 x29|src 302:2  c=2.78961e-19
c3188 x29|src 240:9  c=1.31781e-19
c3187 x29|src 337:2  c=3.14123e-20
c3186 x29|src 353:2  c=4.08423e-20
c3185 x22|src 49:rn  c=6.96726e-19
c3184 x22|src 25:rn  c=6.96726e-19
c3183 x22|src 12:rn  c=1.92142e-19
c3182 x22|src 171:16  c=7.76216e-19
c3181 x22|src 8:rn  c=3.02354e-19
c3180 x22|src 151:16  c=1.30206e-19
cg3179 x16|drn gnd  c=3.84513e-19
c3178 x16|drn 182:16  c=3.74528e-19
c3177 x16|drn 146:16  c=3.7307e-19
c3176 x16|drn 153:16  c=2.32269e-20
c3175 x16|drn 50:rn  c=1.3481e-19
c3174 x16|drn 407:cn  c=9.74156e-21
c3173 x16|drn 188:16  c=4.03631e-19
c3172 x15|src 165:16  c=6.66715e-19
c3171 x15|src 196:q  c=7.76216e-19
c3170 x15|src 145:16  c=6.97923e-19
c3169 x15|src 190:q  c=2.36627e-19
cg3168 530:vdd gnd  c=1.07308e-17
c3167 530:vdd 144:14  c=8.76575e-19
c3166 530:vdd 71:d  c=2.07466e-18
c3165 530:vdd 63:d  c=1.7878e-17
c3164 530:vdd 64:d  c=2.07466e-18
c3163 530:vdd 143:14  c=8.05107e-19
c3162 530:vdd 58:d  c=9.12034e-18
c3161 530:vdd m18|x1|bulk  c=2.7209e-18
c3160 530:vdd 466:gnd  c=5.15371e-21
c3159 530:vdd gnd  c=1.40488e-19
c3158 530:vdd x32|src  c=8.64146e-19
cg3157 529:vdd gnd  c=5.98198e-18
c3156 529:vdd 144:14  c=8.83479e-19
c3155 529:vdd 71:d  c=7.65477e-18
c3154 529:vdd 63:d  c=2.14656e-19
c3153 529:vdd x32|src  c=2.88304e-19
c3152 529:vdd m18|x1|bulk  c=6.97054e-18
c3151 529:vdd 58:d  c=5.88792e-20
c3150 529:vdd 56:d  c=8.69176e-19
cg3149 527:vdd gnd  c=7.64393e-18
c3148 527:vdd 144:14  c=2.83143e-18
c3147 527:vdd 61:d  c=1.12959e-18
c3146 527:vdd 143:14  c=2.88237e-18
c3145 527:vdd x32|src  c=5.11826e-19
c3144 527:vdd m18|x1|bulk  c=6.21869e-18
c3143 527:vdd 56:d  c=1.15858e-18
cg3142 vdd gnd  c=5.25058e-17
c3141 vdd 61:d  c=1.07439e-19
c3140 vdd 144:14  c=5.31184e-17
c3139 vdd 468:gnd  c=8.20252e-21
c3138 vdd 71:d  c=6.2034e-18
c3137 vdd 63:d  c=2.36818e-18
c3136 vdd 64:d  c=3.29311e-18
c3135 vdd 56:d  c=7.08601e-19
c3134 vdd 143:14  c=8.76575e-19
c3133 vdd 32:rn  c=1.70116e-17
c3132 vdd 58:d  c=1.25779e-17
c3131 vdd m18|x1|bulk  c=1.51985e-17
c3130 vdd 466:gnd  c=2.56977e-19
c3129 vdd gnd  c=3.73448e-18
c3128 vdd x32|src  c=2.74519e-19
cg3127 526:vdd gnd  c=6.16141e-18
c3126 526:vdd 66:d  c=2.09514e-19
c3125 526:vdd 65:d  c=7.56186e-18
c3124 526:vdd 135:14  c=1.79434e-18
c3123 526:vdd m18|x1|bulk  c=6.5582e-18
c3122 526:vdd x26|src  c=3.48381e-19
c3121 526:vdd 56:d  c=8.36883e-20
cg3120 525:vdd gnd  c=5.08123e-18
c3119 525:vdd 66:d  c=1.75774e-17
c3118 525:vdd 140:14  c=8.05107e-19
c3117 525:vdd 61:d  c=1.98763e-18
c3116 525:vdd 62:d  c=1.75774e-17
c3115 525:vdd 144:14  c=8.76575e-19
c3114 525:vdd 404:cn  c=7.75046e-21
c3113 525:vdd 331:2  c=1.46422e-21
c3112 525:vdd 56:d  c=2.26394e-17
c3111 525:vdd 143:14  c=8.05107e-19
c3110 525:vdd x26|src  c=8.64146e-19
c3109 525:vdd m18|x1|bulk  c=1.28855e-18
c3108 525:vdd 135:14  c=8.76575e-19
c3107 525:vdd 53:d  c=1.98763e-18
c3106 525:vdd 60:d  c=1.98763e-18
c3105 525:vdd 136:14  c=7.57627e-19
c3104 525:vdd x32|src  c=8.64146e-19
c3103 525:vdd 65:d  c=1.98763e-18
cg3102 523:vdd gnd  c=8.48729e-18
c3101 523:vdd 351:2  c=2.04975e-18
c3100 523:vdd 220:9  c=8.05107e-19
c3099 523:vdd 327:2  c=1.7792e-17
c3098 523:vdd 328:2  c=2.04975e-18
c3097 523:vdd m18|x1|bulk  c=2.76991e-18
c3096 523:vdd x28|drn  c=8.64146e-19
c3095 523:vdd 308:2  c=6.16884e-20
c3094 523:vdd 300:2  c=2.67077e-18
c3093 523:vdd 302:2  c=4.89702e-18
c3092 523:vdd 240:9  c=8.76575e-19
c3091 523:vdd 353:2  c=2.88933e-18
c3090 523:vdd 312:2  c=6.39528e-18
c3089 523:vdd 347:2  c=2.52503e-18
cg3088 522:vdd gnd  c=5.29023e-18
c3087 522:vdd 240:9  c=7.92176e-19
c3086 522:vdd 351:2  c=8.02639e-18
c3085 522:vdd 327:2  c=2.35227e-19
c3084 522:vdd 300:2  c=7.63243e-20
c3083 522:vdd x28|drn  c=2.47303e-19
c3082 522:vdd m18|x1|bulk  c=6.32895e-18
c3081 522:vdd 303:2  c=7.37726e-19
cg3080 520:vdd gnd  c=5.23039e-18
c3079 520:vdd 218:9  c=8.05107e-19
c3078 520:vdd 198:9  c=8.76575e-19
c3077 520:vdd 339:2  c=1.98763e-18
c3076 520:vdd 336:2  c=1.75774e-17
c3075 520:vdd 340:2  c=1.98763e-18
c3074 520:vdd 326:2  c=1.75774e-17
c3073 520:vdd 220:9  c=8.05107e-19
c3072 520:vdd 303:2  c=2.26593e-17
c3071 520:vdd m18|x1|bulk  c=1.43044e-18
c3070 520:vdd x27|src  c=7.76216e-19
c3069 520:vdd x28|drn  c=8.64146e-19
c3068 520:vdd 240:9  c=8.76575e-19
c3067 520:vdd 206:9  c=7.66698e-19
c3066 520:vdd 296:2  c=1.98763e-18
c3065 520:vdd 325:2  c=1.98763e-18
cg3064 519:vdd gnd  c=6.16988e-18
c3063 519:vdd 339:2  c=8.13299e-18
c3062 519:vdd 336:2  c=2.4037e-19
c3061 519:vdd m18|x1|bulk  c=5.8073e-18
c3060 519:vdd 198:9  c=3.86836e-19
c3059 519:vdd 303:2  c=7.33017e-19
cg3058 518:vdd gnd  c=7.21068e-18
c3057 518:vdd 240:9  c=2.93806e-18
c3056 518:vdd 340:2  c=2.88183e-19
c3055 518:vdd 220:9  c=3.61567e-18
c3054 518:vdd m18|x1|bulk  c=5.8073e-18
c3053 518:vdd 303:2  c=1.04321e-18
c3052 518:vdd x28|drn  c=4.6719e-19
cg3051 517:vdd gnd  c=7.78853e-18
c3050 517:vdd 218:9  c=4.94928e-18
c3049 517:vdd m18|x1|bulk  c=5.8073e-18
c3048 517:vdd 198:9  c=3.14879e-18
c3047 517:vdd x27|src  c=3.64552e-19
cg3046 516:vdd gnd  c=7.93317e-18
c3045 516:vdd 435:3  c=4.109e-18
c3044 516:vdd m10|x1|src  c=3.84442e-19
c3043 516:vdd m18|x1|bulk  c=5.8073e-18
c3042 516:vdd 433:3  c=5.58979e-18
c3041 516:vdd 206:9  c=7.81442e-20
cg3040 514:vdd gnd  c=6.67909e-18
c3039 514:vdd 230:9  c=2.15257e-17
c3038 514:vdd m10|x1|gate  c=6.85142e-18
c3037 514:vdd m10|x1|src  c=7.77302e-19
c3036 514:vdd m11|x1|drn  c=8.67977e-19
c3035 514:vdd m18|x1|bulk  c=3.28586e-18
c3034 514:vdd 434:3  c=9.61062e-19
c3033 514:vdd 51:rn  c=9.52594e-19
c3032 514:vdd 431:3  c=8.05107e-19
c3031 514:vdd 237:9  c=4.71428e-19
c3030 514:vdd 435:3  c=9.31789e-19
c3029 514:vdd 40:rn  c=1.98268e-18
c3028 514:vdd 433:3  c=8.05107e-19
c3027 514:vdd 27:rn  c=1.75508e-17
c3026 514:vdd 43:rn  c=7.32044e-18
c3025 514:vdd 44:rn  c=1.96335e-19
cg3024 513:vdd gnd  c=7.25554e-18
c3023 513:vdd m11|x1|drn  c=3.67035e-19
c3022 513:vdd m11|x1|gate  c=2.11584e-18
c3021 513:vdd 354:cn  c=6.76249e-18
c3020 513:vdd 338:2  c=2.00761e-19
c3019 513:vdd 310:2  c=1.5245e-19
c3018 513:vdd m18|x1|bulk  c=5.8073e-18
c3017 513:vdd 434:3  c=2.6255e-18
c3016 513:vdd 370:cn  c=3.02532e-21
cg3015 512:vdd gnd  c=6.33659e-18
c3014 512:vdd 435:3  c=3.42942e-19
c3013 512:vdd 237:9  c=2.17848e-20
c3012 512:vdd 232:9  c=6.58004e-20
c3011 512:vdd 230:9  c=6.71507e-18
c3010 512:vdd m18|x1|bulk  c=6.32909e-18
c3009 512:vdd m10|x1|gate  c=2.09412e-18
cg3008 511:vdd gnd  c=7.96208e-18
c3007 511:vdd 338:2  c=3.22569e-18
c3006 511:vdd 322:2  c=5.61097e-18
c3005 511:vdd 370:cn  c=1.88781e-21
c3004 511:vdd m18|x1|bulk  c=5.8073e-18
c3003 511:vdd m11|x1|src  c=3.82304e-19
cg3002 510:vdd gnd  c=7.81753e-18
c3001 510:vdd 239:9  c=3.18369e-18
c3000 510:vdd x12|src  c=3.63093e-19
c2999 510:vdd m18|x1|bulk  c=5.8073e-18
c2998 510:vdd 216:9  c=4.94928e-18
cg2997 509:vdd gnd  c=5.88217e-18
c2996 509:vdd x11|drn  c=2.45091e-19
c2995 509:vdd 367:cn  c=8.43058e-19
c2994 509:vdd 293:4  c=2.15513e-18
c2993 509:vdd 239:9  c=1.98398e-19
c2992 509:vdd 392:cn  c=8.07523e-18
c2991 509:vdd m18|x1|bulk  c=5.8073e-18
c2990 509:vdd 393:cn  c=2.35227e-19
cg2989 508:vdd gnd  c=7.21833e-18
c2988 508:vdd 293:4  c=3.39491e-18
c2987 508:vdd 390:cn  c=2.87226e-19
c2986 508:vdd 269:4  c=3.59389e-18
c2985 508:vdd m18|x1|bulk  c=5.8073e-18
c2984 508:vdd 367:cn  c=1.17557e-18
c2983 508:vdd x11|drn  c=4.64792e-19
cg2982 507:vdd gnd  c=7.18991e-18
c2981 507:vdd 390:cn  c=7.78304e-20
c2980 507:vdd 367:cn  c=1.13094e-18
c2979 507:vdd 208:9  c=3.79618e-18
c2978 507:vdd 202:9  c=2.78826e-18
c2977 507:vdd x10|drn  c=4.5346e-19
c2976 507:vdd m18|x1|bulk  c=5.8073e-18
cg2975 506:vdd gnd  c=6.12736e-18
c2974 506:vdd x10|drn  c=2.3473e-19
c2973 506:vdd 412:cn  c=8.16843e-18
c2972 506:vdd 289:4  c=5.46647e-19
c2971 506:vdd 202:9  c=6.28976e-19
c2970 506:vdd 389:cn  c=2.4037e-19
c2969 506:vdd 367:cn  c=7.91669e-19
c2968 506:vdd 368:cn  c=7.69386e-21
c2967 506:vdd m18|x1|bulk  c=5.8073e-18
cg2966 505:vdd gnd  c=7.83303e-18
c2965 505:vdd 289:4  c=4.029e-18
c2964 505:vdd 252:4  c=4.92338e-18
c2963 505:vdd x10|src  c=3.64863e-19
c2962 505:vdd m18|x1|bulk  c=5.8073e-18
cg2961 503:vdd gnd  c=1.16704e-17
c2960 503:vdd 25:rn  c=2.04873e-18
c2959 503:vdd x21|src  c=8.64146e-19
c2958 503:vdd 48:rn  c=2.89432e-18
c2957 503:vdd 6:rn  c=2.79741e-18
c2956 503:vdd 8:rn  c=5.58759e-18
c2955 503:vdd 412:cn  c=2.73439e-20
c2954 503:vdd 289:4  c=2.63542e-18
c2953 503:vdd 171:16  c=8.05107e-19
c2952 503:vdd 389:cn  c=2.43562e-19
c2951 503:vdd 367:cn  c=2.73439e-20
c2950 503:vdd 158:16  c=2.69348e-21
c2949 503:vdd 151:16  c=8.76575e-19
c2948 503:vdd 252:4  c=6.57679e-18
c2947 503:vdd 49:rn  c=2.04873e-18
c2946 503:vdd 26:rn  c=1.77884e-17
cg2945 501:vdd gnd  c=7.81535e-18
c2944 501:vdd 184:16  c=5.19807e-23
c2943 501:vdd 147:16  c=3.15816e-18
c2942 501:vdd 169:16  c=4.93511e-18
c2941 501:vdd 247:4  c=3.07546e-19
c2940 501:vdd x19|src  c=3.56622e-19
c2939 501:vdd m18|x1|bulk  c=5.8073e-18
cg2938 500:vdd gnd  c=7.149e-18
c2937 500:vdd 4:rn  c=2.23485e-17
c2936 500:vdd x21|src  c=8.64146e-19
c2935 500:vdd 171:16  c=8.05107e-19
c2934 500:vdd 3:rn  c=1.98763e-18
c2933 500:vdd 22:rn  c=1.98763e-18
c2932 500:vdd 147:16  c=8.76575e-19
c2931 500:vdd 151:16  c=8.76575e-19
c2930 500:vdd 33:rn  c=1.98763e-18
c2929 500:vdd 34:rn  c=1.75774e-17
c2928 500:vdd 23:rn  c=1.98763e-18
c2927 500:vdd 24:rn  c=1.75774e-17
c2926 500:vdd 247:4  c=7.14629e-19
c2925 500:vdd 157:16  c=7.51194e-19
c2924 500:vdd x19|src  c=8.64146e-19
c2923 500:vdd 169:16  c=8.05107e-19
cg2922 498:vdd gnd  c=6.51034e-18
c2921 498:vdd 281:4  c=2.22698e-17
c2920 498:vdd 266:4  c=1.98763e-18
c2919 498:vdd 267:4  c=1.75774e-17
c2918 498:vdd 245:4  c=1.98763e-18
c2917 498:vdd 147:16  c=8.76575e-19
c2916 498:vdd 292:4  c=1.98763e-18
c2915 498:vdd 167:16  c=8.05107e-19
c2914 498:vdd 268:4  c=1.75774e-17
c2913 498:vdd 276:4  c=1.98763e-18
c2912 498:vdd x17|drn  c=8.64146e-19
c2911 498:vdd 247:4  c=7.14629e-19
c2910 498:vdd 157:16  c=1.62777e-18
c2909 498:vdd x19|src  c=8.64146e-19
c2908 498:vdd 169:16  c=8.05107e-19
cg2907 497:vdd gnd  c=7.50508e-18
c2906 497:vdd 281:4  c=1.15362e-18
c2905 497:vdd 266:4  c=2.88183e-19
c2904 497:vdd 157:16  c=2.93089e-18
c2903 497:vdd x17|drn  c=4.64639e-19
c2902 497:vdd m18|x1|bulk  c=5.8073e-18
c2901 497:vdd 167:16  c=3.61314e-18
cg2900 495:vdd gnd  c=6.50896e-18
c2899 495:vdd 281:4  c=7.78429e-19
c2898 495:vdd 278:4  c=8.02639e-18
c2897 495:vdd 263:4  c=2.35227e-19
c2896 495:vdd 157:16  c=7.86498e-19
c2895 495:vdd x17|drn  c=2.45053e-19
c2894 495:vdd m18|x1|bulk  c=5.8073e-18
cg2893 494:vdd gnd  c=5.82368e-18
c2892 494:vdd 292:4  c=8.13299e-18
c2891 494:vdd 281:4  c=7.70781e-19
c2890 494:vdd 268:4  c=2.4037e-19
c2889 494:vdd m18|x1|bulk  c=5.8073e-18
c2888 494:vdd 147:16  c=3.86836e-19
cg2887 492:vdd gnd  c=1.45075e-17
c2886 492:vdd x9|drn  c=4.53294e-19
c2885 492:vdd m18|x1|bulk  c=5.8073e-18
c2884 492:vdd 249:4  c=2.77778e-19
cg2883 491:vdd gnd  c=7.88102e-18
c2882 491:vdd 261:4  c=5.61097e-18
c2881 491:vdd 153:16  c=1.91916e-20
c2880 491:vdd 249:4  c=3.24438e-18
c2879 491:vdd x9|src  c=3.82998e-19
c2878 491:vdd m18|x1|bulk  c=5.8073e-18
cg2877 489:vdd gnd  c=1.38528e-17
c2876 489:vdd 190:q  c=8.76575e-19
c2875 489:vdd 261:4  c=6.35179e-18
c2874 489:vdd 145:16  c=2.07323e-18
c2873 489:vdd x14|drn  c=8.64146e-19
c2872 489:vdd 441:gnd  c=1.58687e-19
c2871 489:vdd 153:16  c=5.05071e-19
c2870 489:vdd 249:4  c=2.53131e-18
c2869 489:vdd 165:16  c=2.05008e-18
c2868 489:vdd 166:16  c=1.77931e-17
c2867 489:vdd 196:q  c=8.05107e-19
cg2866 488:vdd gnd  c=6.24281e-18
c2865 488:vdd 166:16  c=2.35227e-19
c2864 488:vdd 165:16  c=8.0264e-18
c2863 488:vdd 153:16  c=1.27808e-20
c2862 488:vdd 152:16  c=8.26483e-19
c2861 488:vdd m18|x1|bulk  c=5.98582e-18
c2860 488:vdd x14|drn  c=2.45053e-19
c2859 488:vdd 190:q  c=7.86897e-19
cg2858 486:vdd gnd  c=6.59852e-18
c2857 486:vdd 189:q  c=1.61864e-18
c2856 486:vdd 190:q  c=8.76575e-19
c2855 486:vdd 148:16  c=1.98763e-18
c2854 486:vdd 192:q  c=8.05107e-19
c2853 486:vdd x13|src  c=7.76216e-19
c2852 486:vdd x14|drn  c=8.64146e-19
c2851 486:vdd 159:16  c=1.98763e-18
c2850 486:vdd 160:16  c=1.75774e-17
c2849 486:vdd 152:16  c=2.48008e-17
c2848 486:vdd 153:16  c=1.01429e-20
c2847 486:vdd 163:16  c=1.98763e-18
c2846 486:vdd 164:16  c=1.75774e-17
c2845 486:vdd 196:q  c=8.05107e-19
cg2844 484:vdd gnd  c=6.61719e-18
c2843 484:vdd 160:16  c=2.4037e-19
c2842 484:vdd 159:16  c=8.133e-18
c2841 484:vdd m18|x1|bulk  c=6.42015e-18
c2840 484:vdd 152:16  c=7.71809e-19
c2839 484:vdd 189:q  c=3.87026e-19
cg2838 483:vdd gnd  c=7.60371e-18
c2837 483:vdd 163:16  c=2.88183e-19
c2836 483:vdd 196:q  c=3.61314e-18
c2835 483:vdd m18|x1|bulk  c=6.05112e-18
c2834 483:vdd 152:16  c=1.15662e-18
c2833 483:vdd 190:q  c=2.9316e-18
c2832 483:vdd x14|drn  c=4.64639e-19
cg2831 482:vdd gnd  c=1.00571e-17
c2830 482:vdd 193:q  c=1.5694e-21
c2829 482:vdd 192:q  c=4.94928e-18
c2828 482:vdd m18|x1|bulk  c=9.89449e-18
c2827 482:vdd 189:q  c=3.14928e-18
c2826 482:vdd x13|src  c=3.64552e-19
cg2825 481:vdd gnd  c=1.08394e-17
c2824 481:vdd 181:16  c=1.82982e-19
c2823 481:vdd 182:16  c=2.9627e-19
c2822 481:vdd 279:4  c=5.04161e-18
c2821 481:vdd 278:4  c=2.05008e-18
c2820 481:vdd 263:4  c=1.77931e-17
c2819 481:vdd 281:4  c=2.07323e-18
c2818 481:vdd 146:16  c=1.39119e-19
c2817 481:vdd 167:16  c=8.05107e-19
c2816 481:vdd x17|drn  c=8.64146e-19
c2815 481:vdd 290:4  c=2.89692e-18
c2814 481:vdd 247:4  c=3.37756e-18
c2813 481:vdd 157:16  c=8.76575e-19
c2812 481:vdd 188:16  c=1.52588e-21
c2811 x17|src 290:4  c=1.71931e-19
c2810 x17|src 281:4  c=6.97923e-19
c2809 x17|src 279:4  c=2.5586e-19
c2808 x17|src 278:4  c=6.66715e-19
c2807 x17|src 167:16  c=7.76216e-19
c2806 x17|src 157:16  c=2.36627e-19
cg2805 480:vdd gnd  c=2.02625e-16
c2804 480:vdd 189:q  c=1.56072e-16
c2803 480:vdd 190:q  c=9.93588e-17
c2802 480:vdd 279:4  c=1.61458e-19
c2801 480:vdd 261:4  c=2.6405e-18
c2800 480:vdd 278:4  c=1.15224e-18
c2799 480:vdd 281:4  c=5.60118e-19
c2798 480:vdd 148:16  c=2.84429e-18
c2797 480:vdd 146:16  c=1.26302e-19
c2796 480:vdd 192:q  c=3.49703e-18
c2795 480:vdd x13|src  c=3.33553e-19
c2794 480:vdd x14|drn  c=2.74519e-19
c2793 480:vdd 167:16  c=2.96048e-19
c2792 480:vdd m18|x1|bulk  c=9.84956e-17
c2791 480:vdd 159:16  c=6.36178e-18
c2790 480:vdd 160:16  c=2.36818e-18
c2789 480:vdd 191:q  c=5.37346e-19
c2788 480:vdd 152:16  c=1.34286e-17
c2787 480:vdd 441:gnd  c=8.60372e-19
c2786 480:vdd 153:16  c=4.59761e-19
c2785 480:vdd 50:rn  c=1.08199e-17
c2784 480:vdd x17|drn  c=5.69781e-20
c2783 480:vdd 249:4  c=5.41291e-17
c2782 480:vdd 163:16  c=7.55432e-18
c2781 480:vdd 285:4  c=3.1434e-19
c2780 480:vdd 290:4  c=7.12614e-18
c2779 480:vdd 164:16  c=2.36818e-18
c2778 480:vdd 165:16  c=1.25565e-18
c2777 480:vdd 196:q  c=3.70797e-18
c2776 480:vdd 157:16  c=1.77702e-17
c2775 480:vdd 188:16  c=2.50699e-18
cg2774 479:vdd gnd  c=1.69857e-17
c2773 479:vdd 4:rn  c=9.12339e-18
c2772 479:vdd x21|src  c=2.74519e-19
c2771 479:vdd 289:4  c=1.27843e-19
c2770 479:vdd 171:16  c=8.76575e-19
c2769 479:vdd 3:rn  c=2.84429e-18
c2768 479:vdd 22:rn  c=2.84429e-18
c2767 479:vdd 250:4  c=1.12203e-18
c2766 479:vdd 147:16  c=5.17166e-17
c2765 479:vdd 292:4  c=8.3321e-20
c2764 479:vdd 151:16  c=5.16226e-17
c2763 479:vdd 32:rn  c=5.57418e-18
c2762 479:vdd 33:rn  c=5.71456e-18
c2761 479:vdd 34:rn  c=2.36818e-18
c2760 479:vdd 23:rn  c=5.71456e-18
c2759 479:vdd 24:rn  c=2.36818e-18
c2758 479:vdd 247:4  c=1.75034e-18
c2757 479:vdd 157:16  c=4.70344e-17
c2756 479:vdd x19|src  c=2.74519e-19
c2755 479:vdd 169:16  c=8.76575e-19
c2754 479:vdd 186:16  c=2.09315e-19
c2753 479:vdd 49:rn  c=1.07439e-19
cg2752 478:vdd gnd  c=1.05113e-17
c2751 478:vdd 181:16  c=1.80192e-17
c2750 478:vdd 182:16  c=2.07332e-18
c2749 478:vdd 278:4  c=2.95389e-19
c2748 478:vdd 263:4  c=1.82982e-19
c2747 478:vdd 146:16  c=2.71164e-18
c2746 478:vdd x9|drn  c=5.39429e-19
c2745 478:vdd m18|x1|bulk  c=4.56362e-18
c2744 478:vdd 184:16  c=9.5326e-20
c2743 478:vdd 188:16  c=2.10197e-18
cg2742 477:vdd gnd  c=2.45577e-17
c2741 477:vdd 181:16  c=3.60849e-18
c2740 477:vdd 182:16  c=5.51136e-18
c2739 477:vdd 278:4  c=6.76024e-19
c2738 477:vdd 146:16  c=7.24239e-18
c2737 477:vdd x9|drn  c=1.68959e-19
c2736 477:vdd m18|x1|bulk  c=5.96148e-18
c2735 477:vdd 50:rn  c=1.54944e-17
c2734 477:vdd 249:4  c=3.09242e-17
c2733 477:vdd 157:16  c=3.81281e-18
c2732 477:vdd 188:16  c=5.876e-18
cg2731 476:vdd gnd  c=2.33079e-17
c2730 476:vdd 66:d  c=2.34292e-18
c2729 476:vdd 140:14  c=8.76575e-19
c2728 476:vdd 61:d  c=5.71456e-18
c2727 476:vdd 421:cn  c=2.05897e-19
c2726 476:vdd 144:14  c=5.17866e-17
c2725 476:vdd 62:d  c=2.36818e-18
c2724 476:vdd 350:2  c=8.34767e-20
c2723 476:vdd 71:d  c=1.07439e-19
c2722 476:vdd 319:2  c=9.20859e-19
c2721 476:vdd 307:2  c=1.37373e-18
c2720 476:vdd 56:d  c=9.36764e-18
c2719 476:vdd 143:14  c=8.76575e-19
c2718 476:vdd x26|src  c=1.45971e-19
c2717 476:vdd 32:rn  c=5.60286e-18
c2716 476:vdd m18|x1|bulk  c=8.00702e-18
c2715 476:vdd 135:14  c=5.09543e-17
c2714 476:vdd 53:d  c=2.9983e-18
c2713 476:vdd 60:d  c=2.965e-18
c2712 476:vdd 348:2  c=1.41169e-20
c2711 476:vdd 347:2  c=4.5685e-20
c2710 476:vdd 136:14  c=4.68821e-17
c2709 476:vdd x32|src  c=2.74519e-19
c2708 476:vdd 65:d  c=5.19279e-18
c2707 476:vdd 352:2  c=3.56609e-18
cg2706 475:vdd gnd  c=1.72939e-17
c2705 475:vdd 25:rn  c=3.03004e-18
c2704 475:vdd 4:rn  c=9.16326e-19
c2703 475:vdd x21|src  c=2.74519e-19
c2702 475:vdd 48:rn  c=5.41376e-17
c2701 475:vdd 6:rn  c=2.03284e-18
c2700 475:vdd 8:rn  c=3.67323e-18
c2699 475:vdd 412:cn  c=5.19283e-19
c2698 475:vdd 289:4  c=4.68155e-17
c2697 475:vdd 171:16  c=8.76575e-19
c2696 475:vdd 202:9  c=4.89621e-19
c2695 475:vdd 251:4  c=2.87028e-18
c2694 475:vdd 151:16  c=5.0926e-17
c2693 475:vdd 252:4  c=2.7012e-18
c2692 475:vdd 242:4  c=5.06617e-18
c2691 475:vdd 12:rn  c=1.28109e-17
c2690 475:vdd 23:rn  c=1.07439e-19
c2689 475:vdd 294:4  c=4.82548e-18
c2688 475:vdd 246:4  c=8.31552e-18
c2687 475:vdd 49:rn  c=6.64403e-18
c2686 475:vdd 26:rn  c=2.36818e-18
cg2685 474:vdd gnd  c=2.22727e-17
c2684 474:vdd 278:4  c=1.07439e-19
c2683 474:vdd 281:4  c=1.00097e-17
c2682 474:vdd 266:4  c=5.76916e-18
c2681 474:vdd 267:4  c=2.36818e-18
c2680 474:vdd 245:4  c=2.84429e-18
c2679 474:vdd 147:16  c=5.17028e-17
c2678 474:vdd 292:4  c=5.18199e-18
c2677 474:vdd 32:rn  c=5.57418e-18
c2676 474:vdd 167:16  c=8.76575e-19
c2675 474:vdd 268:4  c=2.36818e-18
c2674 474:vdd 276:4  c=2.84429e-18
c2673 474:vdd m18|x1|bulk  c=5.8073e-18
c2672 474:vdd x17|drn  c=2.74519e-19
c2671 474:vdd 33:rn  c=1.07439e-19
c2670 474:vdd 157:16  c=9.89663e-17
c2669 474:vdd x19|src  c=2.74519e-19
c2668 474:vdd 419:cn  c=1.68543e-19
c2667 474:vdd 169:16  c=8.76575e-19
cg2666 473:vdd gnd  c=4.25163e-17
c2665 473:vdd 190:q  c=5.17853e-17
c2664 473:vdd 261:4  c=2.53131e-18
c2663 473:vdd 145:16  c=3.05606e-18
c2662 473:vdd x14|drn  c=2.74519e-19
c2661 473:vdd m18|x1|bulk  c=6.00394e-18
c2660 473:vdd 152:16  c=9.19894e-19
c2659 473:vdd 153:16  c=3.43745e-18
c2658 473:vdd 50:rn  c=1.94812e-17
c2657 473:vdd 249:4  c=4.77823e-17
c2656 473:vdd 163:16  c=1.07439e-19
c2655 473:vdd 165:16  c=6.08567e-18
c2654 473:vdd 166:16  c=2.36818e-18
c2653 473:vdd 196:q  c=8.76575e-19
cg2652 472:vdd gnd  c=2.0558e-17
c2651 472:vdd 218:9  c=8.76575e-19
c2650 472:vdd 427:3  c=8.0362e-19
c2649 472:vdd 425:3  c=1.34638e-18
c2648 472:vdd 198:9  c=5.09439e-17
c2647 472:vdd 306:2  c=1.95171e-17
c2646 472:vdd 468:gnd  c=2.26196e-20
c2645 472:vdd 339:2  c=5.19976e-18
c2644 472:vdd 336:2  c=2.344e-18
c2643 472:vdd 340:2  c=5.76916e-18
c2642 472:vdd 326:2  c=2.36818e-18
c2641 472:vdd 351:2  c=1.07439e-19
c2640 472:vdd 220:9  c=8.76575e-19
c2639 472:vdd 303:2  c=9.56511e-18
c2638 472:vdd m18|x1|bulk  c=7.43046e-18
c2637 472:vdd x27|src  c=1.30562e-19
c2636 472:vdd x28|drn  c=2.74519e-19
c2635 472:vdd 435:3  c=3.87456e-18
c2634 472:vdd 240:9  c=5.14171e-17
c2633 472:vdd 206:9  c=4.45166e-17
c2632 472:vdd 296:2  c=3.0753e-18
c2631 472:vdd 325:2  c=3.04707e-18
c2630 472:vdd 347:2  c=1.25828e-19
c2629 472:vdd 426:3  c=1.84488e-21
c2628 x31|src 140:14  c=8.64146e-19
c2627 x31|src 61:d  c=5.67946e-19
c2626 x31|src 421:cn  c=1.26562e-19
c2625 x31|src 144:14  c=1.72587e-19
c2624 x31|src 56:d  c=2.99254e-18
c2623 x31|src 363:cn  c=6.73592e-20
c2622 x31|src 143:14  c=8.64146e-19
c2621 x31|src 32:rn  c=1.63619e-19
c2620 x31|src 135:14  c=2.74519e-19
c2619 x31|src 53:d  c=5.67946e-19
c2618 x31|src 60:d  c=5.67946e-19
c2617 x31|src 348:2  c=3.52481e-20
c2616 x31|src 65:d  c=5.67946e-19
cg2615 471:vdd gnd  c=1.73007e-17
c2614 471:vdd 230:9  c=9.18556e-18
c2613 471:vdd 427:3  c=2.77248e-17
c2612 471:vdd 425:3  c=4.89792e-18
c2611 471:vdd 198:9  c=8.91528e-19
c2610 471:vdd 306:2  c=7.56986e-18
c2609 471:vdd m10|x1|gate  c=2.11976e-18
c2608 471:vdd m10|x1|src  c=1.20565e-19
c2607 471:vdd m11|x1|drn  c=1.36078e-19
c2606 471:vdd 338:2  c=1.29001e-18
c2605 471:vdd m18|x1|bulk  c=2.64116e-18
c2604 471:vdd 434:3  c=6.18629e-17
c2603 471:vdd 51:rn  c=1.14654e-17
c2602 471:vdd 431:3  c=7.55128e-19
c2601 471:vdd 237:9  c=1.50375e-17
c2600 471:vdd 435:3  c=5.61774e-17
c2599 471:vdd 206:9  c=5.31156e-19
c2598 471:vdd 40:rn  c=3.97343e-18
c2597 471:vdd 433:3  c=8.10835e-19
c2596 471:vdd 27:rn  c=2.21739e-18
c2595 471:vdd 43:rn  c=7.4621e-18
c2594 471:vdd 45:rn  c=3.80023e-19
c2593 471:vdd 426:3  c=5.2315e-18
cg2592 470:vdd gnd  c=2.33259e-17
c2591 470:vdd 425:3  c=4.22844e-19
c2590 470:vdd 306:2  c=2.0825e-17
c2589 470:vdd 350:2  c=5.09179e-18
c2588 470:vdd 307:2  c=7.84099e-18
c2587 470:vdd 340:2  c=1.07439e-19
c2586 470:vdd 351:2  c=6.11182e-18
c2585 470:vdd 220:9  c=8.76575e-19
c2584 470:vdd 327:2  c=2.36818e-18
c2583 470:vdd 328:2  c=3.33323e-18
c2582 470:vdd 303:2  c=6.11469e-19
c2581 470:vdd m18|x1|bulk  c=6.87552e-18
c2580 470:vdd x28|drn  c=2.74519e-19
c2579 470:vdd 308:2  c=2.5224e-20
c2578 470:vdd 300:2  c=2.15717e-18
c2577 470:vdd 302:2  c=3.94123e-18
c2576 470:vdd 240:9  c=5.11236e-17
c2575 470:vdd 337:2  c=2.85048e-18
c2574 470:vdd 353:2  c=5.21205e-17
c2573 470:vdd 312:2  c=2.85356e-18
c2572 470:vdd 311:2  c=5.27984e-18
c2571 470:vdd 347:2  c=4.40163e-17
c2570 470:vdd 136:14  c=4.81434e-19
cg2569 x27|drn gnd  c=2.70252e-20
c2568 x27|drn 218:9  c=8.64146e-19
c2567 x27|drn 198:9  c=2.74519e-19
c2566 x27|drn 306:2  c=6.02422e-19
c2565 x27|drn 339:2  c=5.67946e-19
c2564 x27|drn 340:2  c=5.67946e-19
c2563 x27|drn 220:9  c=8.64146e-19
c2562 x27|drn 364:cn  c=5.61441e-20
c2561 x27|drn 303:2  c=2.76381e-18
c2560 x27|drn 240:9  c=2.74519e-19
c2559 x27|drn 296:2  c=5.67946e-19
c2558 x27|drn 325:2  c=5.67946e-19
c2557 x23|src 31:rn  c=1.22649e-20
c2556 x23|src 230:9  c=2.78423e-18
c2555 x23|src 200:9  c=7.66172e-20
c2554 x23|src 306:2  c=2.36035e-20
c2553 x23|src 364:cn  c=2.33856e-20
c2552 x23|src 51:rn  c=9.85428e-20
c2551 x23|src 431:3  c=8.63198e-19
c2550 x23|src 433:3  c=8.62964e-19
c2549 x23|src 40:rn  c=5.5746e-19
c2548 x23|src 43:rn  c=1.21351e-18
c2547 x20|src 4:rn  c=3.32368e-18
c2546 x20|src 171:16  c=8.64146e-19
c2545 x20|src 3:rn  c=5.67946e-19
c2544 x20|src 22:rn  c=5.67946e-19
c2543 x20|src 147:16  c=2.74519e-19
c2542 x20|src 151:16  c=2.74519e-19
c2541 x20|src 33:rn  c=5.67946e-19
c2540 x20|src 23:rn  c=5.67946e-19
c2539 x20|src 169:16  c=8.64146e-19
c2538 x18|drn 281:4  c=3.02023e-18
c2537 x18|drn 266:4  c=5.67946e-19
c2536 x18|drn 245:4  c=5.67946e-19
c2535 x18|drn 147:16  c=2.74519e-19
c2534 x18|drn 292:4  c=5.67946e-19
c2533 x18|drn 167:16  c=8.64146e-19
c2532 x18|drn 276:4  c=5.67946e-19
c2531 x18|drn 157:16  c=2.74519e-19
c2530 x18|drn 169:16  c=8.64146e-19
cg2529 469:vdd gnd  c=2.24245e-17
c2528 469:vdd 182:16  c=5.4461e-19
c2527 469:vdd 279:4  c=3.99565e-18
c2526 469:vdd 278:4  c=6.08567e-18
c2525 469:vdd 263:4  c=2.36818e-18
c2524 469:vdd 281:4  c=3.82894e-18
c2523 469:vdd 266:4  c=1.07439e-19
c2522 469:vdd 167:16  c=8.76575e-19
c2521 469:vdd m18|x1|bulk  c=5.8073e-18
c2520 469:vdd 50:rn  c=6.69332e-18
c2519 469:vdd x17|drn  c=2.74519e-19
c2518 469:vdd 249:4  c=3.83311e-18
c2517 469:vdd 285:4  c=2.15212e-18
c2516 469:vdd 290:4  c=5.54584e-17
c2515 469:vdd 247:4  c=3.20106e-18
c2514 469:vdd 157:16  c=5.07115e-17
c2513 469:vdd 188:16  c=4.25854e-19
c2512 x13|drn 163:16  c=5.67946e-19
c2511 x13|drn 196:q  c=8.64146e-19
c2510 x13|drn 159:16  c=5.67946e-19
c2509 x13|drn 192:q  c=8.64146e-19
c2508 x13|drn 152:16  c=3.58582e-18
c2507 x13|drn 190:q  c=2.74519e-19
c2506 x13|drn 148:16  c=5.67946e-19
c2505 x13|drn 189:q  c=2.74519e-19
cg2504 m11|x1|bulk gnd  c=1.86549e-16
c2503 m11|x1|bulk 340:2  c=1.52797e-17
c2502 m11|x1|bulk 326:2  c=3.83169e-18
c2501 m11|x1|bulk 351:2  c=1.45691e-17
c2500 m11|x1|bulk 327:2  c=4.07148e-18
c2499 m11|x1|bulk 328:2  c=8.67947e-18
c2498 m11|x1|bulk 303:2  c=5.39872e-17
c2497 m11|x1|bulk 433:3  c=8.96592e-18
c2496 m11|x1|bulk 145:16  c=7.24303e-18
c2495 m11|x1|bulk 148:16  c=6.70968e-18
c2494 m11|x1|bulk 459:gnd  c=7.98612e-20
c2493 m11|x1|bulk 146:16  c=8.41341e-18
c2492 m11|x1|bulk 308:2  c=6.15765e-19
c2491 m11|x1|bulk 302:2  c=5.85966e-18
c2490 m11|x1|bulk 218:9  c=1.16145e-17
c2489 m11|x1|bulk 147:16  c=7.39268e-18
c2488 m11|x1|bulk 151:16  c=5.96659e-18
c2487 m11|x1|bulk 65:d  c=1.34464e-17
c2486 m11|x1|bulk 66:d  c=3.83169e-18
c2485 m11|x1|bulk 135:14  c=6.73375e-18
c2484 m11|x1|bulk 220:9  c=7.15617e-18
c2483 m11|x1|bulk 61:d  c=1.48487e-17
c2482 m11|x1|bulk 62:d  c=3.83169e-18
c2481 m11|x1|bulk 53:d  c=7.56968e-18
c2480 m11|x1|bulk 221:9  c=1.40559e-19
c2479 m11|x1|bulk 60:d  c=7.56968e-18
c2478 m11|x1|bulk 404:cn  c=4.97532e-19
c2477 m11|x1|bulk 54:d  c=5.89328e-18
c2476 m11|x1|bulk 71:d  c=1.49826e-17
c2475 m11|x1|bulk 63:d  c=4.08603e-18
c2474 m11|x1|bulk 64:d  c=8.44541e-18
c2473 m11|x1|bulk 56:d  c=5.40809e-17
c2472 m11|x1|bulk 462:gnd  c=1.51243e-19
c2471 m11|x1|bulk 58:d  c=5.8532e-18
c2470 m11|x1|bulk 59:d  c=6.63955e-18
c2469 m11|x1|bulk 437:gnd  c=3.3502e-19
c2468 m11|x1|bulk 436:gnd  c=2.29201e-19
c2467 m11|x1|bulk 438:gnd  c=2.64252e-19
c2466 m11|x1|bulk 138:14  c=8.25247e-18
c2465 m11|x1|bulk 439:gnd  c=2.71107e-19
c2464 m11|x1|bulk 441:gnd  c=3.4829e-19
c2463 m11|x1|bulk 329:2  c=8.21293e-18
c2462 m11|x1|bulk 249:4  c=1.06555e-17
c2461 m11|x1|bulk 140:14  c=1.09825e-17
c2460 m11|x1|bulk 290:4  c=2.38005e-18
c2459 m11|x1|bulk 157:16  c=7.77874e-18
c2458 m11|x1|bulk 331:2  c=1.17995e-19
c2457 m11|x1|bulk 419:cn  c=6.05391e-19
c2456 m11|x1|bulk 186:16  c=1.84347e-18
c2455 m11|x1|bulk 143:14  c=7.37774e-18
c2454 m11|x1|bulk 142:14  c=1.40565e-19
c2453 m11|x1|bulk 48:rn  c=1.80427e-18
c2452 m11|x1|bulk 289:4  c=1.87589e-18
c2451 m11|x1|bulk 418:cn  c=5.97675e-19
c2450 m11|x1|bulk 202:9  c=4.01701e-18
c2449 m11|x1|bulk 466:gnd  c=1.60165e-19
c2448 m11|x1|bulk 251:4  c=8.64812e-19
c2447 m11|x1|bulk 189:q  c=1.29527e-17
c2446 m11|x1|bulk 239:9  c=7.59744e-18
c2445 m11|x1|bulk 190:q  c=6.8342e-18
c2444 m11|x1|bulk 420:cn  c=1.35669e-19
c2443 m11|x1|bulk 338:2  c=6.43035e-18
c2442 m11|x1|bulk 310:2  c=6.61473e-19
c2441 m11|x1|bulk 434:3  c=2.13499e-18
c2440 m11|x1|bulk 51:rn  c=7.45099e-19
c2439 m11|x1|bulk 237:9  c=9.28756e-19
c2438 m11|x1|bulk 356:cn  c=7.23271e-18
c2437 m11|x1|bulk 359:cn  c=6.70063e-18
c2436 m11|x1|bulk 435:3  c=2.65804e-18
c2435 m11|x1|bulk 238:9  c=6.05359e-19
c2434 m11|x1|bulk 240:9  c=5.27905e-18
c2433 m11|x1|bulk 354:cn  c=3.70222e-17
c2432 m11|x1|bulk 206:9  c=6.28222e-20
c2431 m11|x1|bulk 337:2  c=4.99967e-19
c2430 m11|x1|bulk 353:2  c=1.42104e-18
c2429 m11|x1|bulk 311:2  c=3.89017e-18
c2428 m11|x1|bulk 348:2  c=2.17149e-18
c2427 m11|x1|bulk 347:2  c=2.68872e-18
c2426 m11|x1|bulk 136:14  c=4.48645e-18
c2425 m11|x1|bulk 352:2  c=1.25869e-18
c2424 m11|x1|bulk 421:cn  c=1.02054e-18
c2423 m11|x1|bulk 144:14  c=5.75131e-18
c2422 m11|x1|bulk 72:d  c=7.79329e-18
c2421 m11|x1|bulk 422:cn  c=3.08549e-19
c2420 m11|x1|bulk 252:4  c=1.14106e-17
c2419 m11|x1|bulk 3:rn  c=6.70968e-18
c2418 m11|x1|bulk 22:rn  c=6.70968e-18
c2417 m11|x1|bulk 2:rn  c=6.84558e-18
c2416 m11|x1|bulk 312:2  c=1.29523e-17
c2415 m11|x1|bulk 50:rn  c=7.8607e-18
c2414 m11|x1|bulk 407:cn  c=1.08548e-18
c2413 m11|x1|bulk 362:cn  c=4.36223e-19
c2412 m11|x1|bulk 12:rn  c=5.72673e-18
c2411 m11|x1|bulk 294:4  c=4.46707e-18
c2410 m11|x1|bulk 355:cn  c=2.78794e-19
c2409 m11|x1|bulk 259:4  c=4.87636e-18
c2408 m11|x1|bulk 246:4  c=3.82755e-18
c2407 m11|x1|bulk 192:q  c=1.36089e-17
c2406 m11|x1|bulk 426:3  c=4.91735e-18
c2405 m11|x1|bulk 31:rn  c=1.00002e-18
c2404 m11|x1|bulk 193:q  c=1.8894e-20
c2403 m11|x1|bulk 427:3  c=2.59646e-18
c2402 m11|x1|bulk 425:3  c=4.69802e-18
c2401 m11|x1|bulk 212:9  c=4.50158e-19
c2400 m11|x1|bulk 200:9  c=1.33063e-18
c2399 m11|x1|bulk 306:2  c=1.39769e-17
c2398 m11|x1|bulk 350:2  c=4.24587e-18
c2397 m11|x1|bulk gnd  c=4.08671e-19
c2396 m11|x1|bulk 319:2  c=5.3119e-18
c2395 m11|x1|bulk 445:gnd  c=1.6308e-20
c2394 m11|x1|bulk 307:2  c=4.03323e-18
c2393 m11|x1|bulk 363:cn  c=7.24782e-19
c2392 m11|x1|bulk 20:rn  c=2.47811e-18
c2391 m11|x1|bulk 32:rn  c=1.60569e-17
c2390 m11|x1|bulk 364:cn  c=4.43625e-18
c2389 m11|x1|bulk 196:q  c=7.11363e-18
c2388 m11|x1|bulk 159:16  c=1.51587e-17
c2387 m11|x1|bulk 152:16  c=6.88876e-17
c2386 m11|x1|bulk 153:16  c=1.06106e-17
c2385 m11|x1|bulk m10|x1|gate  c=5.70417e-19
c2384 m11|x1|bulk 163:16  c=1.52797e-17
c2383 m11|x1|bulk 261:4  c=1.12846e-17
c2382 m11|x1|bulk 165:16  c=1.4586e-17
c2381 m11|x1|bulk m11|x1|gate  c=5.73876e-19
c2380 m11|x1|bulk 188:16  c=1.0739e-17
c2379 m11|x1|bulk 182:16  c=1.98465e-17
c2378 m11|x1|bulk 279:4  c=1.11264e-17
c2377 m11|x1|bulk 167:16  c=7.11363e-18
c2376 m11|x1|bulk 278:4  c=1.4586e-17
c2375 m11|x1|bulk 281:4  c=6.22962e-17
c2374 m11|x1|bulk 266:4  c=1.52797e-17
c2373 m11|x1|bulk 365:cn  c=4.2723e-19
c2372 m11|x1|bulk 396:cn  c=7.68331e-20
c2371 m11|x1|bulk 292:4  c=1.34483e-17
c2370 m11|x1|bulk 276:4  c=6.70968e-18
c2369 m11|x1|bulk 169:16  c=8.29049e-18
c2368 m11|x1|bulk 184:16  c=2.51817e-19
c2367 m11|x1|bulk 33:rn  c=1.5481e-17
c2366 m11|x1|bulk 442:gnd  c=1.98635e-20
c2365 m11|x1|bulk 23:rn  c=1.5481e-17
c2364 m11|x1|bulk 440:gnd  c=2.07326e-20
c2363 m11|x1|bulk 247:4  c=1.86348e-17
c2362 m11|x1|bulk 171:16  c=8.20706e-18
c2361 m11|x1|bulk 49:rn  c=1.65935e-17
c2360 m11|x1|bulk 158:16  c=2.04242e-20
c2359 m11|x1|bulk 25:rn  c=7.23766e-18
c2358 m11|x1|bulk 4:rn  c=5.66591e-17
c2357 m11|x1|bulk 8:rn  c=7.30614e-18
c2356 m11|x1|bulk 412:cn  c=1.45758e-17
c2355 m11|x1|bulk 367:cn  c=6.82551e-17
c2354 m11|x1|bulk 368:cn  c=7.05296e-18
c2353 m11|x1|bulk 208:9  c=7.06078e-18
c2352 m11|x1|bulk 390:cn  c=1.52916e-17
c2351 m11|x1|bulk 392:cn  c=1.46023e-17
c2350 m11|x1|bulk 198:9  c=7.02577e-18
c2349 m11|x1|bulk 269:4  c=7.07719e-18
c2348 m11|x1|bulk 370:cn  c=2.07477e-19
c2347 m11|x1|bulk 245:4  c=6.70968e-18
c2346 m11|x1|bulk 243:4  c=6.21271e-18
c2345 m11|x1|bulk 215:9  c=8.78695e-21
c2344 m11|x1|bulk 216:9  c=1.15276e-17
c2343 m11|x1|bulk 40:rn  c=1.12161e-17
c2342 m11|x1|bulk 242:4  c=2.93629e-18
c2341 m11|x1|bulk 43:rn  c=2.39713e-17
c2340 m11|x1|bulk 322:2  c=1.13405e-17
c2339 m11|x1|bulk 230:9  c=3.61085e-17
c2338 m11|x1|bulk 203:9  c=1.74702e-18
c2337 m11|x1|bulk 296:2  c=7.99968e-18
c2336 m11|x1|bulk 325:2  c=8.68115e-18
c2335 m11|x1|bulk 232:9  c=2.8653e-18
c2334 m11|x1|bulk 297:2  c=6.72198e-18
c2333 m11|x1|bulk 321:2  c=1.37417e-19
c2332 m11|x1|bulk 234:9  c=1.08099e-19
c2331 m11|x1|bulk 339:2  c=1.46014e-17
c2330 m11|x1|bulk 431:3  c=1.08548e-17
c2329 m11|x1|bulk 336:2  c=4.07541e-18
cg2328 468:gnd gnd  c=5.07964e-16
c2327 468:gnd 418:cn  c=1.84347e-17
c2326 468:gnd 355:cn  c=1.06511e-17
c2325 468:gnd 185:16  c=2.43051e-18
c2324 468:gnd m7|x1|drn  c=2.44244e-19
c2323 468:gnd 250:4  c=4.94347e-18
c2322 468:gnd 251:4  c=6.61395e-19
c2321 468:gnd 303:2  c=4.15493e-19
c2320 468:gnd 291:4  c=3.10382e-18
c2319 468:gnd x1|drn  c=1.12929e-19
c2318 468:gnd x1|src  c=1.09871e-20
c2317 468:gnd 205:9  c=1.18379e-18
c2316 468:gnd 235:9  c=5.65302e-17
c2315 468:gnd 131:c  c=3.39987e-19
c2314 468:gnd 342:2  c=1.02922e-18
c2313 468:gnd 405:cn  c=2.74647e-18
c2312 468:gnd 420:cn  c=1.32779e-17
c2311 468:gnd 349:2  c=4.55802e-17
c2310 468:gnd x4|src  c=5.46084e-19
c2309 468:gnd 51:rn  c=3.41245e-18
c2308 468:gnd 212:9  c=1.51919e-17
c2307 468:gnd 284:4  c=1.68846e-18
c2306 468:gnd x5|drn  c=3.09951e-19
c2305 468:gnd 200:9  c=8.46205e-17
c2304 468:gnd 158:16  c=2.52777e-18
c2303 468:gnd 4:rn  c=8.39254e-20
c2302 468:gnd 238:9  c=6.33268e-17
c2301 468:gnd 206:9  c=3.74135e-18
c2300 468:gnd 37:rn  c=2.21167e-18
c2299 468:gnd 207:9  c=4.93043e-17
c2298 468:gnd 126:c  c=2.49971e-19
c2297 468:gnd 363:cn  c=3.13538e-18
c2296 468:gnd 353:2  c=2.37884e-20
c2295 468:gnd 82:c  c=3.0544e-18
c2294 468:gnd 311:2  c=9.27131e-19
c2293 468:gnd 348:2  c=2.56887e-16
c2292 468:gnd 368:cn  c=1.41836e-18
c2291 468:gnd 136:14  c=1.69609e-19
c2290 468:gnd 364:cn  c=6.53724e-17
c2289 468:gnd 221:9  c=2.63855e-18
c2288 468:gnd 404:cn  c=1.67965e-19
c2287 468:gnd 133:c  c=3.31198e-19
c2286 468:gnd 394:cn  c=2.71184e-18
c2285 468:gnd 421:cn  c=3.1638e-18
c2284 468:gnd 198:9  c=8.58151e-21
c2283 468:gnd 137:14  c=5.33447e-17
c2282 468:gnd 56:d  c=2.55241e-20
c2281 468:gnd 270:4  c=4.69638e-17
c2280 468:gnd x2|src  c=6.30175e-20
c2279 468:gnd 69:d  c=1.02922e-18
c2278 468:gnd 87:c  c=4.45559e-17
c2277 468:gnd 249:4  c=7.75466e-17
c2276 468:gnd 43:rn  c=1.51595e-21
c2275 468:gnd 45:rn  c=3.07388e-19
c2274 468:gnd 157:16  c=4.77058e-20
c2273 468:gnd 39:rn  c=4.17416e-18
c2272 468:gnd 331:2  c=3.65542e-18
c2271 468:gnd 419:cn  c=6.07961e-18
c2270 468:gnd 203:9  c=2.21975e-18
c2269 468:gnd 186:16  c=1.40956e-17
c2268 468:gnd 156:16  c=1.12866e-20
c2267 468:gnd 396:cn  c=1.69297e-19
c2266 468:gnd 231:9  c=2.43981e-18
c2265 468:gnd 264:4  c=2.70347e-18
c2264 468:gnd 295:4  c=3.75733e-19
c2263 468:gnd 388:cn  c=2.37945e-18
c2262 468:gnd 234:9  c=5.10435e-18
c2261 468:gnd 142:14  c=3.57155e-18
c2260 468:gnd 187:16  c=4.54027e-17
c2259 468:gnd m5|x1|drn  c=4.74677e-20
c2258 468:gnd 407:cn  c=2.62059e-18
c2257 468:gnd 362:cn  c=5.71896e-18
c2256 x8|drn 69:d  c=7.43977e-19
c2255 x8|drn 32:rn  c=1.1177e-19
c2254 x8|drn 137:14  c=5.22628e-19
c2253 x8|drn 82:c  c=2.59898e-20
c2252 x8|drn 57:d  c=7.43977e-19
c2251 x8|drn 142:14  c=7.76216e-19
c2250 x8|drn 58:d  c=2.50354e-19
c2249 x8|drn 364:cn  c=1.04564e-19
c2248 m5|x1|src 306:2  c=9.42699e-20
c2247 m5|x1|src 82:c  c=9.62429e-22
c2246 m5|x1|src 32:rn  c=1.2035e-19
c2245 m5|x1|src 221:9  c=7.76216e-19
c2244 m5|x1|src 364:cn  c=2.93215e-19
c2243 m5|x1|src 341:2  c=7.01546e-19
c2242 m5|x1|src 345:2  c=4.18252e-20
c2241 m5|x1|src 342:2  c=7.43977e-19
c2240 m5|x1|src 308:2  c=2.63096e-19
c2239 m5|x1|src 302:2  c=9.25333e-20
c2238 m5|x1|src 207:9  c=5.31818e-19
c2237 m5|x1|src 353:2  c=5.96693e-20
c2236 m5|x1|src 311:2  c=3.4663e-19
c2235 m5|x1|src 348:2  c=5.68768e-19
cg2234 x7|drn gnd  c=5.0469e-20
c2233 x7|drn 39:rn  c=1.0201e-19
c2232 x7|drn 203:9  c=1.38125e-18
c2231 x7|drn 212:9  c=2.72628e-19
c2230 x7|drn 204:9  c=3.79516e-19
c2229 x7|drn 231:9  c=3.72738e-19
c2228 x7|drn 232:9  c=1.07858e-19
c2227 x7|drn 305:2  c=1.02329e-19
c2226 x7|drn 233:9  c=8.61539e-20
c2225 x7|drn 234:9  c=1.35604e-18
c2224 x7|drn 82:c  c=7.27244e-20
c2223 x7|drn 32:rn  c=8.94679e-20
c2222 x7|drn 364:cn  c=6.02166e-20
c2221 x7|drn 238:9  c=1.85813e-19
c2220 x7|drn 104:c  c=1.17376e-19
c2219 x7|drn 206:9  c=2.65506e-19
c2218 x7|drn 41:rn  c=1.0201e-19
c2217 x3|src 37:rn  c=5.37911e-20
c2216 x3|src 409:cn  c=1.85005e-19
c2215 x3|src 388:cn  c=1.85005e-19
c2214 x3|src 82:c  c=7.37235e-20
c2213 x3|src 32:rn  c=6.06054e-20
c2212 x3|src 364:cn  c=4.35007e-19
c2211 x3|src 155:16  c=3.68609e-19
c2210 x3|src 185:16  c=3.9841e-19
c2209 x3|src 183:16  c=7.7319e-20
c2208 x3|src 249:4  c=2.62506e-19
c2207 x3|src 247:4  c=1.8373e-19
c2206 x3|src 157:16  c=5.33498e-20
c2205 x3|src 284:4  c=1.75675e-19
c2204 x3|src 186:16  c=3.14638e-19
c2203 m23|x1|src 162:16  c=7.43977e-19
c2202 m23|x1|src 191:q  c=4.82322e-19
c2201 m23|x1|src 154:16  c=7.40118e-19
c2200 m23|x1|src 193:q  c=7.76216e-19
c2199 m23|x1|src 189:q  c=2.30414e-19
c2198 m23|x1|src 153:16  c=1.07328e-18
cg2197 466:gnd gnd  c=1.12663e-17
c2196 466:gnd 137:14  c=8.76575e-19
c2195 466:gnd 57:d  c=1.99526e-17
c2194 466:gnd 142:14  c=8.05107e-19
c2193 466:gnd 69:d  c=2.07466e-18
c2192 466:gnd 58:d  c=3.29817e-19
c2191 466:gnd x2|drn  c=8.64146e-19
cg2190 gnd gnd  c=4.24926e-17
c2189 gnd 137:14  c=5.3384e-17
c2188 gnd 57:d  c=6.33236e-18
c2187 gnd 82:c  c=1.45291e-18
c2186 gnd 142:14  c=8.76575e-19
c2185 gnd 69:d  c=4.18643e-18
c2184 gnd 58:d  c=1.87166e-18
c2183 gnd 364:cn  c=2.12943e-17
c2182 gnd x2|drn  c=5.69709e-19
c2181 gnd 348:2  c=3.75126e-18
cg2180 465:gnd gnd  c=8.38815e-18
c2179 465:gnd 69:d  c=6.57207e-18
c2178 465:gnd 137:14  c=1.87116e-18
c2177 465:gnd 58:d  c=8.55331e-21
c2176 465:gnd 57:d  c=2.3604e-19
c2175 465:gnd 56:d  c=5.02694e-23
cg2174 463:gnd gnd  c=7.79888e-18
c2173 463:gnd 346:2  c=2.08577e-19
c2172 463:gnd 342:2  c=6.19166e-18
c2171 463:gnd 207:9  c=7.19384e-19
c2170 463:gnd 311:2  c=3.1423e-20
c2169 463:gnd 308:2  c=4.78566e-20
cg2168 462:gnd gnd  c=6.07524e-18
c2167 462:gnd 331:2  c=6.18556e-20
c2166 462:gnd 221:9  c=8.05107e-19
c2165 462:gnd 341:2  c=1.74897e-18
c2164 462:gnd 345:2  c=3.26884e-19
c2163 462:gnd 346:2  c=1.7878e-17
c2162 462:gnd 342:2  c=2.07466e-18
c2161 462:gnd 308:2  c=4.07994e-19
c2160 462:gnd 302:2  c=8.80829e-20
c2159 462:gnd 207:9  c=8.76575e-19
c2158 462:gnd m5|x1|drn  c=7.76216e-19
c2157 462:gnd 311:2  c=1.07455e-18
c2156 462:gnd 348:2  c=5.47419e-18
cg2155 461:gnd gnd  c=9.06674e-18
c2154 461:gnd 221:9  c=5.61097e-18
c2153 461:gnd 207:9  c=3.19931e-18
c2152 461:gnd 303:2  c=2.92243e-21
c2151 461:gnd m5|x1|drn  c=3.84155e-19
cg2150 459:gnd gnd  c=5.44923e-18
c2149 459:gnd 46:rn  c=1.04103e-18
c2148 459:gnd 39:rn  c=1.84868e-19
c2147 459:gnd 203:9  c=1.18454e-17
c2146 459:gnd 204:9  c=2.00995e-17
c2145 459:gnd 231:9  c=2.07487e-18
c2144 459:gnd 232:9  c=3.32489e-21
c2143 459:gnd x6|src  c=5.39429e-19
c2142 459:gnd 234:9  c=6.30529e-18
c2141 459:gnd 238:9  c=2.30189e-18
c2140 459:gnd 206:9  c=1.71622e-19
c2139 459:gnd 41:rn  c=1.84868e-19
cg2138 458:gnd gnd  c=1.09131e-17
c2137 458:gnd 51:rn  c=2.48699e-19
c2136 458:gnd 349:2  c=2.24163e-19
c2135 458:gnd 45:rn  c=8.71546e-20
c2134 458:gnd 43:rn  c=7.01811e-21
c2133 458:gnd m7|x1|drn  c=4.58366e-19
c2132 458:gnd 87:c  c=1.09884e-17
cg2131 457:gnd gnd  c=9.05071e-18
c2130 457:gnd 77:c  c=4.02554e-19
c2129 457:gnd 87:c  c=2.09504e-17
c2128 457:gnd m7|x1|src  c=1.91313e-19
cg2127 456:gnd gnd  c=8.21629e-18
c2126 456:gnd x1|src  c=1.91313e-19
c2125 456:gnd 77:c  c=4.02554e-19
c2124 456:gnd 87:c  c=2.09251e-17
cg2123 455:gnd gnd  c=7.14959e-18
c2122 455:gnd 77:c  c=3.39989e-19
c2121 455:gnd 87:c  c=1.58254e-17
cg2120 454:gnd gnd  c=8.5754e-18
c2119 454:gnd 270:4  c=8.72514e-18
c2118 454:gnd 367:cn  c=2.39406e-20
c2117 454:gnd x1|drn  c=3.84155e-19
cg2116 453:gnd gnd  c=7.59548e-18
c2115 453:gnd 187:16  c=3.18428e-18
c2114 453:gnd x5|drn  c=1.18308e-18
c2113 453:gnd 158:16  c=4.54218e-18
c2112 453:gnd 8:rn  c=3.45204e-20
c2111 453:gnd 6:rn  c=2.46523e-21
cg2110 452:gnd gnd  c=7.88339e-18
c2109 452:gnd 187:16  c=3.54551e-19
c2108 452:gnd 186:16  c=3.86092e-19
c2107 452:gnd 37:rn  c=6.46791e-18
c2106 452:gnd x4|src  c=8.59994e-19
c2105 452:gnd 5:rn  c=2.07071e-19
c2104 x4|drn 295:4  c=3.92548e-19
c2103 x4|drn 186:16  c=3.15517e-19
c2102 x4|drn 32:rn  c=1.80399e-19
c2101 x4|drn 157:16  c=5.4395e-20
c2100 x4|drn 247:4  c=1.61402e-19
c2099 x4|drn 364:cn  c=6.10353e-19
cg2098 449:gnd gnd  c=8.82898e-18
c2097 449:gnd 419:cn  c=5.20755e-19
c2096 449:gnd 410:cn  c=2.07071e-19
c2095 449:gnd 184:16  c=3.46561e-20
c2094 449:gnd 183:16  c=3.98458e-21
c2093 449:gnd 388:cn  c=6.29887e-18
c2092 449:gnd 249:4  c=2.62744e-19
c2091 449:gnd 146:16  c=3.25053e-21
cg2090 448:gnd gnd  c=8.53518e-18
c2089 448:gnd 184:16  c=3.15539e-20
c2088 448:gnd 396:cn  c=1.91561e-20
c2087 448:gnd 264:4  c=5.60671e-18
c2086 448:gnd 249:4  c=2.78509e-18
c2085 448:gnd 146:16  c=1.54145e-21
c2084 448:gnd m18|x1|src  c=3.8303e-19
cg2083 446:gnd gnd  c=8.05585e-18
c2082 446:gnd 162:16  c=6.19166e-18
c2081 446:gnd 161:16  c=2.08577e-19
c2080 446:gnd 153:16  c=2.07098e-19
c2079 446:gnd 191:q  c=7.19384e-19
cg2078 445:gnd gnd  c=6.84803e-18
c2077 445:gnd 189:q  c=2.30272e-19
c2076 445:gnd 193:q  c=8.05107e-19
c2075 445:gnd 191:q  c=8.76575e-19
c2074 445:gnd 152:16  c=6.93573e-21
c2073 445:gnd 153:16  c=4.70618e-18
c2072 445:gnd 154:16  c=2.08225e-18
c2071 445:gnd 249:4  c=1.9242e-18
c2070 445:gnd m23|x1|drn  c=7.76216e-19
c2069 445:gnd 161:16  c=1.7878e-17
c2068 445:gnd 162:16  c=2.07466e-18
cg2067 443:gnd gnd  c=1.02209e-17
c2066 443:gnd 193:q  c=5.61097e-18
c2065 443:gnd 192:q  c=1.70738e-21
c2064 443:gnd 191:q  c=3.19931e-18
c2063 443:gnd m23|x1|drn  c=3.84155e-19
cg2062 442:gnd gnd  c=1.03215e-17
c2061 442:gnd 4:rn  c=4.16663e-21
c2060 442:gnd 5:rn  c=1.96292e-20
c2059 442:gnd 409:cn  c=7.38131e-20
c2058 442:gnd 410:cn  c=6.57481e-19
c2057 442:gnd 388:cn  c=7.38131e-20
c2056 442:gnd m18|x1|drn  c=5.39429e-19
c2055 442:gnd 155:16  c=2.00926e-17
c2054 442:gnd 185:16  c=2.10374e-18
c2053 442:gnd 183:16  c=1.97246e-21
c2052 442:gnd 247:4  c=2.14249e-19
c2051 442:gnd 157:16  c=1.5699e-20
c2050 442:gnd 288:4  c=8.82602e-19
c2049 442:gnd 284:4  c=2.42083e-19
c2048 442:gnd 186:16  c=3.27641e-18
cg2047 441:gnd gnd  c=2.37025e-16
c2046 441:gnd 189:q  c=1.4593e-17
c2045 441:gnd 190:q  c=3.8271e-19
c2044 441:gnd 193:q  c=3.52814e-18
c2043 441:gnd 388:cn  c=9.27779e-20
c2042 441:gnd 241:4  c=4.07906e-18
c2041 441:gnd 191:q  c=1.11831e-16
c2040 441:gnd 152:16  c=7.12415e-20
c2039 441:gnd 277:4  c=1.44909e-17
c2038 441:gnd 153:16  c=2.86055e-17
c2037 441:gnd 118:c  c=3.89595e-18
c2036 441:gnd 184:16  c=6.3025e-20
c2035 441:gnd 154:16  c=3.96248e-18
c2034 441:gnd 407:cn  c=3.46303e-17
c2033 441:gnd 161:16  c=2.36818e-18
c2032 441:gnd 249:4  c=2.1893e-16
c2031 441:gnd m23|x1|drn  c=3.44141e-19
c2030 441:gnd 162:16  c=5.18891e-18
c2029 441:gnd 264:4  c=2.08632e-19
c2028 441:gnd 132:c  c=2.35853e-19
c2027 441:gnd 157:16  c=2.26603e-20
cg2026 440:gnd gnd  c=1.01576e-17
c2025 440:gnd 4:rn  c=3.26833e-21
c2024 440:gnd 295:4  c=2.8005e-19
c2023 440:gnd x4|src  c=5.57673e-19
c2022 440:gnd 5:rn  c=8.05107e-19
c2021 440:gnd 409:cn  c=1.76859e-20
c2020 440:gnd 155:16  c=1.01575e-18
c2019 440:gnd 247:4  c=1.05539e-19
c2018 440:gnd 287:4  c=2.61662e-19
c2017 440:gnd 288:4  c=2.21759e-17
c2016 440:gnd 186:16  c=3.4294e-18
cg2015 439:gnd gnd  c=8.65494e-18
c2014 439:gnd 187:16  c=3.12804e-18
c2013 439:gnd 365:cn  c=2.59305e-19
c2012 439:gnd 409:cn  c=8.14958e-19
c2011 439:gnd 410:cn  c=8.14958e-19
c2010 439:gnd 388:cn  c=8.14958e-19
c2009 439:gnd 241:4  c=5.4094e-19
c2008 439:gnd 364:cn  c=1.51567e-17
c2007 439:gnd m18|x1|drn  c=9.3469e-20
c2006 439:gnd 277:4  c=1.37848e-18
c2005 439:gnd 155:16  c=9.03038e-18
c2004 439:gnd 185:16  c=5.88538e-18
c2003 439:gnd 249:4  c=2.7325e-17
c2002 439:gnd 285:4  c=2.59538e-19
c2001 439:gnd 247:4  c=1.01575e-20
c2000 439:gnd 157:16  c=4.7423e-20
c1999 439:gnd 288:4  c=1.01324e-19
c1998 439:gnd 284:4  c=6.04184e-19
c1997 439:gnd 186:16  c=3.88197e-17
c1996 439:gnd 156:16  c=3.77309e-20
cg1995 438:gnd gnd  c=9.22103e-18
c1994 438:gnd 295:4  c=1.68505e-18
c1993 438:gnd x4|src  c=2.96099e-19
c1992 438:gnd 5:rn  c=2.40484e-18
c1991 438:gnd 37:rn  c=9.39269e-19
c1990 438:gnd 187:16  c=3.43237e-17
c1989 438:gnd 365:cn  c=4.04806e-19
c1988 438:gnd 251:4  c=4.04892e-19
c1987 438:gnd 291:4  c=2.02516e-19
c1986 438:gnd 364:cn  c=1.557e-17
c1985 438:gnd 277:4  c=6.83129e-19
c1984 438:gnd 155:16  c=1.61322e-18
c1983 438:gnd 185:16  c=4.36715e-19
c1982 438:gnd 249:4  c=3.16705e-18
c1981 438:gnd 285:4  c=2.6041e-19
c1980 438:gnd 87:c  c=5.68428e-19
c1979 438:gnd 157:16  c=2.10659e-20
c1978 438:gnd 287:4  c=1.5649e-19
c1977 438:gnd 286:4  c=2.55029e-18
c1976 438:gnd 270:4  c=8.85049e-19
c1975 438:gnd 288:4  c=1.00905e-17
c1974 438:gnd 284:4  c=7.01023e-18
c1973 438:gnd 186:16  c=4.47361e-17
cg1972 437:gnd gnd  c=1.7761e-17
c1971 437:gnd 212:9  c=1.49741e-18
c1970 437:gnd 200:9  c=5.92529e-19
c1969 437:gnd 331:2  c=2.70224e-19
c1968 437:gnd 394:cn  c=6.64354e-20
c1967 437:gnd 82:c  c=2.82106e-18
c1966 437:gnd 221:9  c=8.76575e-19
c1965 437:gnd 364:cn  c=2.35841e-17
c1964 437:gnd 341:2  c=3.83379e-18
c1963 437:gnd 345:2  c=1.06504e-19
c1962 437:gnd 346:2  c=2.34765e-18
c1961 437:gnd 342:2  c=4.16414e-18
c1960 437:gnd 308:2  c=1.34715e-18
c1959 437:gnd 302:2  c=3.05567e-20
c1958 437:gnd 238:9  c=9.87758e-19
c1957 437:gnd 207:9  c=5.29006e-17
c1956 437:gnd 337:2  c=1.57975e-19
c1955 437:gnd m5|x1|drn  c=3.285e-19
c1954 437:gnd 311:2  c=8.96017e-18
c1953 437:gnd 348:2  c=4.98618e-17
cg1952 m18|x1|bulk gnd  c=2.46245e-17
c1951 m18|x1|bulk 303:2  c=4.07887e-17
c1950 m18|x1|bulk 341:2  c=1.42547e-16
c1949 m18|x1|bulk 345:2  c=1.96743e-19
c1948 m18|x1|bulk 342:2  c=1.45948e-17
c1947 m18|x1|bulk 146:16  c=6.27945e-17
c1946 m18|x1|bulk 308:2  c=9.49936e-17
c1945 m18|x1|bulk 149:16  c=9.49669e-17
c1944 m18|x1|bulk 300:2  c=3.02546e-17
c1943 m18|x1|bulk 302:2  c=3.05447e-17
c1942 m18|x1|bulk 218:9  c=4.66235e-18
c1941 m18|x1|bulk 147:16  c=1.56931e-18
c1940 m18|x1|bulk 128:c  c=4.08082e-17
c1939 m18|x1|bulk 151:16  c=9.64143e-19
c1938 m18|x1|bulk 88:c  c=1.0615e-16
c1937 m18|x1|bulk 126:c  c=5.86398e-17
c1936 m18|x1|bulk 135:14  c=1.90861e-18
c1935 m18|x1|bulk 220:9  c=1.29415e-18
c1934 m18|x1|bulk 221:9  c=1.9139e-17
c1933 m18|x1|bulk 404:cn  c=6.50157e-17
c1932 m18|x1|bulk 54:d  c=1.85004e-18
c1931 m18|x1|bulk 403:cn  c=4.99411e-17
c1930 m18|x1|bulk 394:cn  c=1.62303e-17
c1929 m18|x1|bulk 56:d  c=3.79981e-17
c1928 m18|x1|bulk 57:d  c=2.03337e-16
c1927 m18|x1|bulk 69:d  c=1.33316e-17
c1926 m18|x1|bulk 58:d  c=6.14599e-17
c1925 m18|x1|bulk 59:d  c=4.00103e-17
c1924 m18|x1|bulk 191:q  c=1.29796e-16
c1923 m18|x1|bulk 138:14  c=1.43674e-18
c1922 m18|x1|bulk 329:2  c=1.4234e-18
c1921 m18|x1|bulk 249:4  c=1.54648e-16
c1920 m18|x1|bulk 140:14  c=4.69937e-18
c1919 m18|x1|bulk 132:c  c=9.24453e-18
c1918 m18|x1|bulk 285:4  c=5.58774e-17
c1917 m18|x1|bulk 290:4  c=8.21928e-18
c1916 m18|x1|bulk 157:16  c=3.22231e-17
c1915 m18|x1|bulk 331:2  c=2.0851e-17
c1914 m18|x1|bulk 419:cn  c=1.37613e-17
c1913 m18|x1|bulk 186:16  c=5.72441e-17
c1912 m18|x1|bulk 156:16  c=9.66091e-18
c1911 m18|x1|bulk 143:14  c=1.29415e-18
c1910 m18|x1|bulk 295:4  c=6.84552e-18
c1909 m18|x1|bulk 142:14  c=1.4673e-17
c1908 m18|x1|bulk 187:16  c=1.83841e-17
c1907 m18|x1|bulk 48:rn  c=6.70597e-18
c1906 m18|x1|bulk 289:4  c=1.00129e-18
c1905 m18|x1|bulk 418:cn  c=2.25139e-17
c1904 m18|x1|bulk 202:9  c=1.81191e-17
c1903 m18|x1|bulk 250:4  c=5.56946e-17
c1902 m18|x1|bulk 251:4  c=2.62497e-17
c1901 m18|x1|bulk 291:4  c=1.79923e-18
c1900 m18|x1|bulk 189:q  c=4.48114e-17
c1899 m18|x1|bulk 239:9  c=2.24597e-18
c1898 m18|x1|bulk 190:q  c=3.44058e-18
c1897 m18|x1|bulk 205:9  c=2.11155e-17
c1896 m18|x1|bulk 235:9  c=5.61055e-19
c1895 m18|x1|bulk 131:c  c=7.25601e-18
c1894 m18|x1|bulk 420:cn  c=7.79119e-18
c1893 m18|x1|bulk 338:2  c=6.5943e-19
c1892 m18|x1|bulk 310:2  c=9.36486e-18
c1891 m18|x1|bulk 349:2  c=3.01258e-17
c1890 m18|x1|bulk 51:rn  c=9.47387e-18
c1889 m18|x1|bulk 237:9  c=1.56923e-18
c1888 m18|x1|bulk 238:9  c=2.04071e-17
c1887 m18|x1|bulk 240:9  c=8.21074e-19
c1886 m18|x1|bulk 354:cn  c=1.28403e-16
c1885 m18|x1|bulk 206:9  c=6.22205e-17
c1884 m18|x1|bulk 207:9  c=3.48497e-17
c1883 m18|x1|bulk 337:2  c=5.82505e-19
c1882 m18|x1|bulk 353:2  c=7.76428e-18
c1881 m18|x1|bulk 311:2  c=3.82824e-17
c1880 m18|x1|bulk 348:2  c=1.44996e-16
c1879 m18|x1|bulk 347:2  c=1.53164e-18
c1878 m18|x1|bulk 136:14  c=5.80618e-17
c1877 m18|x1|bulk 352:2  c=6.47674e-19
c1876 m18|x1|bulk 133:c  c=2.84706e-17
c1875 m18|x1|bulk 421:cn  c=1.31779e-17
c1874 m18|x1|bulk 144:14  c=1.69893e-18
c1873 m18|x1|bulk 75:c  c=4.60323e-17
c1872 m18|x1|bulk 137:14  c=2.75252e-17
c1871 m18|x1|bulk 77:c  c=3.56534e-17
c1870 m18|x1|bulk 89:c  c=9.26451e-17
c1869 m18|x1|bulk 72:d  c=2.91469e-17
c1868 m18|x1|bulk 134:c  c=2.30288e-17
c1867 m18|x1|bulk 52:rn  c=1.96051e-17
c1866 m18|x1|bulk 422:cn  c=3.92972e-17
c1865 m18|x1|bulk 2:rn  c=7.38286e-18
c1864 m18|x1|bulk 76:c  c=9.24836e-18
c1863 m18|x1|bulk 312:2  c=4.58619e-18
c1862 m18|x1|bulk 277:4  c=3.15171e-18
c1861 m18|x1|bulk 118:c  c=2.32136e-17
c1860 m18|x1|bulk 50:rn  c=3.49178e-17
c1859 m18|x1|bulk 407:cn  c=4.1399e-17
c1858 m18|x1|bulk 362:cn  c=6.03851e-18
c1857 m18|x1|bulk 1:rn  c=2.21744e-18
c1856 m18|x1|bulk 12:rn  c=5.8799e-18
c1855 m18|x1|bulk 355:cn  c=1.33585e-17
c1854 m18|x1|bulk 259:4  c=3.14922e-18
c1853 m18|x1|bulk 246:4  c=3.86721e-18
c1852 m18|x1|bulk 236:9  c=3.0671e-18
c1851 m18|x1|bulk 81:c  c=1.03039e-17
c1850 m18|x1|bulk 405:cn  c=7.16652e-18
c1849 m18|x1|bulk 304:2  c=4.29217e-18
c1848 m18|x1|bulk 31:rn  c=2.40709e-18
c1847 m18|x1|bulk 193:q  c=2.07862e-17
c1846 m18|x1|bulk 212:9  c=1.64674e-17
c1845 m18|x1|bulk 200:9  c=4.36341e-17
c1844 m18|x1|bulk 305:2  c=2.03992e-17
c1843 m18|x1|bulk 306:2  c=1.18299e-17
c1842 m18|x1|bulk 319:2  c=4.33829e-18
c1841 m18|x1|bulk 307:2  c=6.15781e-18
c1840 m18|x1|bulk 74:c  c=1.01222e-17
c1839 m18|x1|bulk 363:cn  c=1.23916e-17
c1838 m18|x1|bulk 82:c  c=5.7197e-17
c1837 m18|x1|bulk 83:c  c=1.00072e-17
c1836 m18|x1|bulk 20:rn  c=1.47089e-17
c1835 m18|x1|bulk 32:rn  c=8.29349e-17
c1834 m18|x1|bulk 364:cn  c=1.06343e-16
c1833 m18|x1|bulk 387:cn  c=1.59379e-17
c1832 m18|x1|bulk 152:16  c=4.0123e-17
c1831 m18|x1|bulk 153:16  c=4.6679e-16
c1830 m18|x1|bulk 154:16  c=6.28673e-17
c1829 m18|x1|bulk 162:16  c=1.55528e-17
c1828 m18|x1|bulk 261:4  c=4.52499e-18
c1827 m18|x1|bulk 103:c  c=8.15341e-17
c1826 m18|x1|bulk 111:c  c=1.0249e-17
c1825 m18|x1|bulk 182:16  c=3.10103e-17
c1824 m18|x1|bulk 279:4  c=1.54261e-17
c1823 m18|x1|bulk 281:4  c=1.39255e-17
c1822 m18|x1|bulk 365:cn  c=5.3035e-17
c1821 m18|x1|bulk 396:cn  c=2.46926e-17
c1820 m18|x1|bulk 264:4  c=2.01657e-17
c1819 m18|x1|bulk 409:cn  c=8.66009e-18
c1818 m18|x1|bulk 388:cn  c=1.1116e-17
c1817 m18|x1|bulk 155:16  c=1.28319e-16
c1816 m18|x1|bulk 185:16  c=1.3437e-17
c1815 m18|x1|bulk 184:16  c=1.36224e-16
c1814 m18|x1|bulk 183:16  c=3.59603e-17
c1813 m18|x1|bulk 247:4  c=1.61764e-16
c1812 m18|x1|bulk 283:4  c=1.71317e-17
c1811 m18|x1|bulk 287:4  c=3.94309e-17
c1810 m18|x1|bulk 286:4  c=9.55679e-17
c1809 m18|x1|bulk 284:4  c=1.49322e-17
c1808 m18|x1|bulk 158:16  c=2.07636e-17
c1807 m18|x1|bulk 4:rn  c=1.78666e-17
c1806 m18|x1|bulk 5:rn  c=1.42655e-16
c1805 m18|x1|bulk 37:rn  c=1.38545e-17
c1804 m18|x1|bulk 6:rn  c=2.87645e-17
c1803 m18|x1|bulk 8:rn  c=2.84685e-17
c1802 m18|x1|bulk 367:cn  c=4.16962e-17
c1801 m18|x1|bulk 368:cn  c=2.00969e-16
c1800 m18|x1|bulk 120:c  c=8.57961e-18
c1799 m18|x1|bulk 121:c  c=1.02913e-17
c1798 m18|x1|bulk 198:9  c=2.06193e-18
c1797 m18|x1|bulk 270:4  c=2.65692e-17
c1796 m18|x1|bulk 123:c  c=2.46583e-18
c1795 m18|x1|bulk 84:c  c=7.12401e-17
c1794 m18|x1|bulk 86:c  c=3.51778e-17
c1793 m18|x1|bulk 370:cn  c=6.98036e-17
c1792 m18|x1|bulk 243:4  c=1.13293e-17
c1791 m18|x1|bulk 104:c  c=1.45221e-17
c1790 m18|x1|bulk 215:9  c=1.34521e-17
c1789 m18|x1|bulk 87:c  c=1.02861e-16
c1788 m18|x1|bulk 241:4  c=5.45568e-18
c1787 m18|x1|bulk 242:4  c=1.3469e-18
c1786 m18|x1|bulk 43:rn  c=2.18646e-17
c1785 m18|x1|bulk 44:rn  c=1.82693e-17
c1784 m18|x1|bulk 45:rn  c=3.54197e-17
c1783 m18|x1|bulk 41:rn  c=1.00905e-16
c1782 m18|x1|bulk 39:rn  c=9.83265e-18
c1781 m18|x1|bulk 322:2  c=4.22742e-18
c1780 m18|x1|bulk 230:9  c=5.34147e-18
c1779 m18|x1|bulk 203:9  c=1.99096e-16
c1778 m18|x1|bulk 204:9  c=1.81239e-17
c1777 m18|x1|bulk 231:9  c=1.23939e-17
c1776 m18|x1|bulk 232:9  c=3.91033e-17
c1775 m18|x1|bulk 297:2  c=1.0724e-17
c1774 m18|x1|bulk 321:2  c=1.6428e-17
c1773 m18|x1|bulk 233:9  c=2.5982e-17
c1772 m18|x1|bulk 234:9  c=4.66169e-17
cg1771 436:gnd gnd  c=1.89126e-17
c1770 436:gnd 46:rn  c=1.52182e-18
c1769 436:gnd 39:rn  c=1.52182e-18
c1768 436:gnd 203:9  c=1.37185e-17
c1767 436:gnd 212:9  c=7.25789e-18
c1766 436:gnd 200:9  c=4.77669e-17
c1765 436:gnd 204:9  c=9.42329e-18
c1764 436:gnd 231:9  c=6.07772e-18
c1763 436:gnd 233:9  c=8.14452e-19
c1762 436:gnd 234:9  c=4.0165e-18
c1761 436:gnd x6|src  c=7.26759e-20
c1760 436:gnd 82:c  c=3.92545e-18
c1759 436:gnd 235:9  c=5.16034e-20
c1758 436:gnd 364:cn  c=1.31861e-17
c1757 436:gnd 349:2  c=1.22342e-17
c1756 436:gnd 342:2  c=2.16447e-20
c1755 436:gnd 238:9  c=4.0372e-17
c1754 436:gnd 206:9  c=3.85778e-18
c1753 436:gnd 207:9  c=1.62472e-19
c1752 436:gnd 87:c  c=2.26002e-18
c1751 436:gnd 41:rn  c=2.00603e-18
cg1750 435:3 gnd  c=4.63801e-18
c1749 435:3 218:9  c=2.72943e-18
c1748 435:3 230:9  c=1.28178e-17
c1747 435:3 203:9  c=1.8415e-19
c1746 435:3 198:9  c=5.11001e-17
c1745 435:3 232:9  c=2.1004e-18
c1744 435:3 306:2  c=4.4145e-18
c1743 435:3 m10|x1|gate  c=2.7991e-19
c1742 435:3 339:2  c=9.86921e-19
c1741 435:3 338:2  c=3.22318e-20
c1740 435:3 237:9  c=3.60703e-17
c1739 435:3 240:9  c=4.24685e-21
c1738 435:3 206:9  c=1.80861e-17
c1737 435:3 325:2  c=6.53355e-19
c1736 435:3 43:rn  c=3.28747e-19
cg1735 434:3 gnd  c=1.55797e-17
c1734 434:3 m7|x1|src  c=3.4306e-20
c1733 434:3 230:9  c=2.7087e-19
c1732 434:3 306:2  c=4.75075e-18
c1731 434:3 239:9  c=2.63142e-18
c1730 434:3 322:2  c=9.35744e-19
c1729 434:3 m11|x1|src  c=1.2847e-19
c1728 434:3 338:2  c=6.14369e-17
c1727 434:3 310:2  c=3.53892e-17
c1726 434:3 349:2  c=1.38886e-18
c1725 434:3 51:rn  c=2.52665e-18
c1724 434:3 40:rn  c=3.89603e-18
c1723 434:3 27:rn  c=2.49984e-18
c1722 434:3 43:rn  c=5.46901e-18
c1721 434:3 45:rn  c=6.24392e-20
cg1720 m10|x1|src gnd  c=1.09944e-19
c1719 m10|x1|src 230:9  c=1.36681e-18
c1718 m10|x1|src 203:9  c=9.00423e-20
c1717 m10|x1|src 200:9  c=4.51695e-20
c1716 m10|x1|src 232:9  c=4.78762e-19
c1715 m10|x1|src 306:2  c=5.92257e-20
c1714 m10|x1|src 237:9  c=1.05611e-19
c1713 m10|x1|src 206:9  c=5.95005e-21
cg1712 433:3 gnd  c=1.42239e-17
c1711 433:3 218:9  c=6.30843e-18
c1710 433:3 230:9  c=1.48243e-17
c1709 433:3 203:9  c=1.49238e-19
c1708 433:3 198:9  c=2.50683e-18
c1707 433:3 232:9  c=2.62441e-18
c1706 433:3 339:2  c=2.95389e-19
c1705 433:3 336:2  c=1.82982e-19
c1704 433:3 237:9  c=2.83231e-18
c1703 433:3 325:2  c=1.52588e-21
cg1702 431:3 gnd  c=2.60193e-17
c1701 431:3 322:2  c=8.05107e-19
c1700 431:3 m11|x1|src  c=7.75182e-19
c1699 431:3 338:2  c=8.02177e-19
c1698 431:3 310:2  c=3.42918e-18
c1697 431:3 321:2  c=6.84427e-20
c1696 431:3 40:rn  c=1.98736e-18
c1695 431:3 27:rn  c=1.75612e-17
c1694 431:3 43:rn  c=1.98736e-18
cg1693 427:3 gnd  c=2.39376e-17
c1692 427:3 198:9  c=5.39211e-18
c1691 427:3 305:2  c=2.17921e-18
c1690 427:3 306:2  c=4.24556e-17
c1689 427:3 350:2  c=2.56589e-18
c1688 427:3 319:2  c=1.66981e-19
c1687 427:3 307:2  c=3.71652e-18
c1686 427:3 239:9  c=1.25466e-18
c1685 427:3 m11|x1|src  c=1.96912e-19
c1684 427:3 338:2  c=5.27595e-18
cg1683 426:3 gnd  c=3.80515e-17
c1682 426:3 m7|x1|src  c=2.95255e-20
c1681 426:3 305:2  c=3.79964e-18
c1680 426:3 306:2  c=6.39364e-17
c1679 426:3 350:2  c=2.47228e-19
c1678 426:3 307:2  c=1.81785e-19
c1677 426:3 239:9  c=1.54475e-19
c1676 426:3 m11|x1|src  c=4.36485e-20
c1675 426:3 338:2  c=5.21996e-18
c1674 426:3 310:2  c=3.59083e-18
cg1673 425:3 gnd  c=3.08905e-17
c1672 425:3 198:9  c=5.51824e-18
c1671 425:3 305:2  c=3.79964e-18
c1670 425:3 306:2  c=6.48903e-17
c1669 425:3 350:2  c=1.56173e-18
c1668 425:3 319:2  c=4.35603e-20
c1667 425:3 307:2  c=3.61383e-18
c1666 425:3 237:9  c=2.79065e-18
c1665 425:3 206:9  c=1.382e-18
cg1664 m11|x1|drn gnd  c=1.20157e-18
c1663 m11|x1|drn 230:9  c=3.56417e-19
c1662 m11|x1|drn 306:2  c=5.32137e-20
c1661 m11|x1|drn 322:2  c=8.65709e-19
c1660 m11|x1|drn 338:2  c=7.70356e-20
c1659 m11|x1|drn 310:2  c=1.54195e-19
c1658 m11|x1|drn 40:rn  c=5.67734e-19
c1657 m11|x1|drn 43:rn  c=5.67734e-19
cg1656 422:cn gnd  c=3.48752e-17
c1655 422:cn 83:c  c=8.09984e-18
c1654 422:cn 52:rn  c=3.06868e-18
c1653 422:cn 134:c  c=8.63572e-17
c1652 422:cn 137:14  c=1.71399e-17
cg1651 421:cn gnd  c=9.12892e-18
c1650 421:cn 133:c  c=6.64298e-18
c1649 421:cn 137:14  c=9.15519e-17
c1648 421:cn 331:2  c=3.38301e-18
c1647 421:cn 134:c  c=1.29217e-19
c1646 421:cn 74:c  c=7.17966e-19
c1645 421:cn 82:c  c=7.31218e-18
c1644 421:cn 32:rn  c=3.07577e-18
c1643 421:cn 341:2  c=2.69575e-19
c1642 421:cn x2|src  c=3.97549e-19
c1641 421:cn 348:2  c=3.63186e-17
c1640 421:cn 136:14  c=1.18556e-17
cg1639 420:cn gnd  c=5.85204e-18
c1638 420:cn 200:9  c=1.20574e-17
c1637 420:cn 251:4  c=2.20732e-18
c1636 420:cn m11|x1|src  c=2.92117e-20
c1635 420:cn 82:c  c=6.09085e-19
c1634 420:cn 205:9  c=5.3665e-17
c1633 420:cn 131:c  c=7.43588e-17
c1632 420:cn 32:rn  c=4.61469e-19
c1631 420:cn 349:2  c=5.74338e-17
c1630 420:cn 84:c  c=6.03165e-19
c1629 420:cn 86:c  c=4.49162e-18
c1628 420:cn 207:9  c=1.06299e-20
c1627 420:cn 77:c  c=6.65184e-18
c1626 420:cn 89:c  c=1.91631e-18
c1625 420:cn 81:c  c=5.90609e-18
c1624 420:cn 41:rn  c=6.63565e-19
cg1623 419:cn gnd  c=8.52103e-18
c1622 419:cn 5:rn  c=2.72867e-20
c1621 419:cn 187:16  c=6.06575e-19
c1620 419:cn 149:16  c=2.66816e-19
c1619 419:cn 82:c  c=6.43584e-18
c1618 419:cn 32:rn  c=2.4456e-18
c1617 419:cn m18|x1|src  c=3.37208e-19
c1616 419:cn 153:16  c=1.56943e-19
c1615 419:cn 155:16  c=8.19198e-18
c1614 419:cn 118:c  c=8.3888e-19
c1613 419:cn 184:16  c=4.92007e-18
c1612 419:cn 50:rn  c=3.68577e-19
c1611 419:cn 249:4  c=2.95627e-17
c1610 419:cn 264:4  c=3.25604e-18
c1609 419:cn 285:4  c=1.15025e-17
c1608 419:cn 157:16  c=8.94056e-18
c1607 419:cn 286:4  c=2.17132e-19
c1606 419:cn 186:16  c=8.13599e-17
c1605 419:cn 156:16  c=3.05573e-18
cg1604 418:cn gnd  c=1.13847e-17
c1603 418:cn 5:rn  c=2.77667e-18
c1602 418:cn 187:16  c=3.28419e-18
c1601 418:cn 250:4  c=2.51453e-17
c1600 418:cn 251:4  c=3.1534e-17
c1599 418:cn 205:9  c=1.40981e-18
c1598 418:cn 82:c  c=9.21535e-18
c1597 418:cn 32:rn  c=3.02439e-18
c1596 418:cn 89:c  c=1.66864e-18
c1595 418:cn 286:4  c=3.73976e-19
c1594 418:cn 186:16  c=1.81373e-17
cg1593 416:cn gnd  c=5.09855e-19
c1592 416:cn 348:2  c=2.43915e-18
c1591 416:cn 331:2  c=1.7878e-17
c1590 416:cn 142:14  c=1.75794e-17
c1589 416:cn 137:14  c=2.3224e-18
cg1588 412:cn gnd  c=8.17717e-18
c1587 412:cn x10|drn  c=5.60088e-19
c1586 412:cn x10|src  c=6.97848e-19
c1585 412:cn 289:4  c=6.08147e-18
c1584 412:cn 202:9  c=3.38872e-18
c1583 412:cn 293:4  c=1.13472e-19
c1582 412:cn 252:4  c=2.04812e-18
c1581 412:cn 208:9  c=1.98341e-18
c1580 412:cn 23:rn  c=9.11537e-21
c1579 412:cn 49:rn  c=1.10794e-18
c1578 410:cn 249:4  c=3.74864e-18
c1577 410:cn 264:4  c=1.80868e-17
c1576 410:cn 155:16  c=1.38797e-17
cg1575 409:cn gnd  c=1.15848e-18
c1574 409:cn 241:4  c=3.80274e-19
c1573 409:cn m18|x1|src  c=3.64008e-19
c1572 409:cn 155:16  c=1.43021e-17
c1571 409:cn 249:4  c=3.51098e-18
c1570 409:cn 264:4  c=2.09289e-18
c1569 409:cn 285:4  c=2.3619e-20
c1568 409:cn 286:4  c=7.52737e-22
c1567 409:cn 288:4  c=3.48517e-21
cg1566 407:cn gnd  c=4.67352e-17
c1565 407:cn 149:16  c=7.59226e-20
c1564 407:cn 82:c  c=1.86257e-20
c1563 407:cn 241:4  c=1.98972e-18
c1562 407:cn 76:c  c=8.89265e-17
c1561 407:cn 153:16  c=3.21912e-18
c1560 407:cn 277:4  c=5.04987e-17
c1559 407:cn 118:c  c=3.0999e-16
c1558 407:cn 50:rn  c=3.51323e-17
c1557 407:cn 249:4  c=1.04163e-16
c1556 407:cn 132:c  c=7.38212e-18
c1555 407:cn 285:4  c=3.21184e-17
cg1554 405:cn gnd  c=1.13224e-17
c1553 405:cn 349:2  c=7.43992e-18
c1552 405:cn 81:c  c=3.79964e-18
c1551 405:cn 82:c  c=6.57715e-19
c1550 405:cn 205:9  c=5.13751e-18
c1549 405:cn 251:4  c=2.75514e-19
c1548 405:cn 200:9  c=4.68159e-17
cg1547 404:cn gnd  c=1.99952e-17
c1546 404:cn 137:14  c=5.91029e-18
c1545 404:cn 331:2  c=4.01708e-18
c1544 404:cn 348:2  c=3.93752e-18
c1543 404:cn 136:14  c=2.3825e-18
cg1542 403:cn gnd  c=2.15054e-17
c1541 403:cn 348:2  c=4.14514e-18
c1540 403:cn x2|src  c=7.43977e-19
c1539 403:cn x2|drn  c=5.67946e-19
c1538 403:cn 142:14  c=1.98762e-18
c1537 403:cn 331:2  c=2.07466e-18
c1536 403:cn 137:14  c=1.25158e-17
cg1535 396:cn gnd  c=4.93782e-18
c1534 396:cn 146:16  c=7.14726e-21
c1533 396:cn 155:16  c=1.5554e-17
c1532 396:cn 153:16  c=1.28802e-19
c1531 396:cn 184:16  c=2.60134e-19
c1530 396:cn 249:4  c=2.55094e-18
c1529 396:cn 264:4  c=2.50388e-18
c1528 396:cn 285:4  c=1.17806e-18
c1527 396:cn 286:4  c=1.84421e-20
c1526 396:cn 186:16  c=2.01513e-18
c1525 396:cn 156:16  c=1.0728e-19
cg1524 394:cn gnd  c=7.06471e-18
c1523 394:cn 137:14  c=2.93805e-18
c1522 394:cn 331:2  c=2.07466e-18
c1521 394:cn 142:14  c=1.98762e-18
c1520 394:cn x2|drn  c=5.67946e-19
c1519 394:cn x2|src  c=7.43977e-19
c1518 394:cn 348:2  c=3.51055e-18
c1517 393:cn 239:9  c=2.21448e-18
c1516 393:cn 293:4  c=2.48948e-18
c1515 393:cn 269:4  c=1.75618e-17
c1514 393:cn 216:9  c=1.77771e-17
c1513 393:cn 322:2  c=1.82982e-19
cg1512 392:cn gnd  c=8.17888e-18
c1511 392:cn 216:9  c=2.04792e-18
c1510 392:cn x11|drn  c=5.68024e-19
c1509 392:cn x12|src  c=6.57082e-19
c1508 392:cn 293:4  c=5.19691e-18
c1507 392:cn 239:9  c=3.70054e-18
c1506 392:cn 322:2  c=2.94084e-19
c1505 392:cn 338:2  c=6.62482e-19
c1504 392:cn 40:rn  c=5.5013e-21
c1503 392:cn 269:4  c=1.98709e-18
c1502 391:cn 293:4  c=2.46562e-18
c1501 391:cn 208:9  c=1.75547e-17
c1500 391:cn 269:4  c=1.75624e-17
c1499 391:cn 202:9  c=2.2387e-18
cg1498 390:cn gnd  c=8.03828e-18
c1497 390:cn x10|drn  c=5.59444e-19
c1496 390:cn 289:4  c=1.12869e-19
c1495 390:cn x11|drn  c=5.68303e-19
c1494 390:cn 202:9  c=3.37857e-18
c1493 390:cn 293:4  c=4.91835e-18
c1492 390:cn 208:9  c=1.98324e-18
c1491 390:cn 269:4  c=1.98683e-18
c1490 390:cn 49:rn  c=9.11537e-21
c1489 389:cn 289:4  c=2.45865e-18
c1488 389:cn 252:4  c=1.77749e-17
c1487 389:cn 208:9  c=1.75558e-17
c1486 389:cn 202:9  c=2.24715e-18
cg1485 388:cn gnd  c=1.30621e-18
c1484 388:cn m18|x1|src  c=3.64008e-19
c1483 388:cn 185:16  c=1.43021e-17
c1482 388:cn 249:4  c=5.02034e-18
c1481 388:cn 264:4  c=2.09289e-18
c1480 388:cn 284:4  c=1.17653e-20
cg1479 387:cn gnd  c=2.3727e-17
c1478 387:cn 83:c  c=3.79964e-18
c1477 387:cn 137:14  c=3.02664e-18
cg1476 370:cn gnd  c=1.3313e-17
c1475 370:cn 203:9  c=6.02059e-20
c1474 370:cn 322:2  c=1.42585e-19
c1473 370:cn 205:9  c=4.4381e-18
c1472 370:cn m11|x1|src  c=2.87876e-20
c1471 370:cn 131:c  c=5.42492e-18
c1470 370:cn 349:2  c=9.04186e-18
c1469 370:cn 84:c  c=3.24453e-19
c1468 370:cn 86:c  c=1.14509e-17
c1467 370:cn 87:c  c=2.73561e-19
c1466 370:cn 77:c  c=5.93011e-18
c1465 370:cn 89:c  c=4.88219e-18
c1464 370:cn 41:rn  c=3.19424e-18
cg1463 368:cn gnd  c=3.33571e-17
c1462 368:cn 295:4  c=4.41294e-19
c1461 368:cn 5:rn  c=9.48674e-18
c1460 368:cn 48:rn  c=1.9785e-18
c1459 368:cn 6:rn  c=2.61671e-18
c1458 368:cn 8:rn  c=3.40874e-18
c1457 368:cn 202:9  c=1.09829e-17
c1456 368:cn 250:4  c=2.31603e-17
c1455 368:cn 251:4  c=2.02432e-17
c1454 368:cn 2:rn  c=4.2174e-19
c1453 368:cn 239:9  c=3.42849e-19
c1452 368:cn 205:9  c=7.17254e-19
c1451 368:cn 82:c  c=4.25167e-19
c1450 368:cn 310:2  c=9.45091e-20
c1449 368:cn 242:4  c=1.15205e-17
c1448 368:cn 349:2  c=6.07739e-21
c1447 368:cn 84:c  c=1.00732e-18
c1446 368:cn 86:c  c=1.60273e-19
c1445 368:cn 89:c  c=4.10734e-18
c1444 368:cn 283:4  c=1.78646e-20
c1443 368:cn 287:4  c=2.72842e-20
c1442 368:cn 286:4  c=6.85503e-19
c1441 368:cn 43:rn  c=3.8167e-21
c1440 368:cn 45:rn  c=4.86875e-21
c1439 368:cn 186:16  c=3.27437e-18
cg1438 367:cn gnd  c=2.77447e-17
c1437 367:cn 25:rn  c=5.90269e-19
c1436 367:cn 4:rn  c=1.14249e-18
c1435 367:cn x10|drn  c=3.21015e-18
c1434 367:cn x10|src  c=6.97848e-19
c1433 367:cn 289:4  c=4.14266e-18
c1432 367:cn x11|drn  c=3.02728e-18
c1431 367:cn 202:9  c=4.11121e-17
c1430 367:cn 3:rn  c=4.84754e-21
c1429 367:cn 251:4  c=4.55929e-18
c1428 367:cn 293:4  c=1.20762e-17
c1427 367:cn 239:9  c=5.72777e-18
c1426 367:cn 120:c  c=2.2404e-23
c1425 367:cn 252:4  c=2.04812e-18
c1424 367:cn 338:2  c=6.96505e-19
c1423 367:cn 242:4  c=3.97199e-18
c1422 367:cn 123:c  c=3.86387e-22
c1421 367:cn 84:c  c=5.95404e-19
c1420 367:cn 208:9  c=2.456e-17
c1419 367:cn 89:c  c=1.69934e-20
c1418 367:cn 270:4  c=1.12204e-19
c1417 367:cn 43:rn  c=8.09532e-21
c1416 367:cn 269:4  c=2.27608e-17
cg1415 365:cn gnd  c=5.85548e-18
c1414 365:cn 146:16  c=9.97269e-20
c1413 365:cn 149:16  c=1.10571e-19
c1412 365:cn 241:4  c=7.39544e-19
c1411 365:cn 153:16  c=1.27351e-19
c1410 365:cn 155:16  c=4.42995e-17
c1409 365:cn 184:16  c=2.72877e-18
c1408 365:cn 249:4  c=1.1023e-18
c1407 365:cn 264:4  c=8.17887e-20
c1406 365:cn 285:4  c=2.41667e-18
c1405 365:cn 286:4  c=1.78787e-19
c1404 365:cn 186:16  c=2.2909e-18
c1403 365:cn 156:16  c=1.90391e-19
cg1402 364:cn gnd  c=1.16128e-16
c1401 364:cn 250:4  c=7.61783e-18
c1400 364:cn 251:4  c=3.25603e-17
c1399 364:cn 291:4  c=1.50965e-18
c1398 364:cn m7|x1|src  c=1.20744e-19
c1397 364:cn 236:9  c=3.66721e-17
c1396 364:cn 341:2  c=2.12583e-19
c1395 364:cn x1|drn  c=4.29814e-19
c1394 364:cn 205:9  c=2.38052e-17
c1393 364:cn x1|src  c=1.39412e-19
c1392 364:cn 81:c  c=8.88054e-17
c1391 364:cn 235:9  c=1.44459e-18
c1390 364:cn 131:c  c=6.63998e-18
c1389 364:cn 349:2  c=3.67578e-17
c1388 364:cn x4|src  c=2.82235e-19
c1387 364:cn 51:rn  c=4.46896e-18
c1386 364:cn 212:9  c=4.26846e-17
c1385 364:cn x5|drn  c=5.79932e-19
c1384 364:cn 200:9  c=1.12828e-16
c1383 364:cn 238:9  c=8.07457e-18
c1382 364:cn x6|src  c=6.80798e-20
c1381 364:cn 207:9  c=5.12905e-17
c1380 364:cn 74:c  c=9.16053e-17
c1379 364:cn 82:c  c=1.0713e-15
c1378 364:cn 311:2  c=7.3408e-18
c1377 364:cn 83:c  c=8.70805e-17
c1376 364:cn 348:2  c=1.16803e-16
c1375 364:cn 32:rn  c=1.07573e-16
c1374 364:cn 133:c  c=9.21535e-18
c1373 364:cn 137:14  c=3.16594e-17
c1372 364:cn x2|drn  c=2.86548e-19
c1371 364:cn 134:c  c=4.38572e-18
c1370 364:cn 285:4  c=4.08086e-18
c1369 364:cn m11|x1|src  c=3.91386e-20
c1368 364:cn x24|drn  c=5.61441e-20
c1367 364:cn 41:rn  c=4.25167e-19
c1366 364:cn 203:9  c=1.00647e-18
c1365 364:cn x26|src  c=1.04871e-20
c1364 364:cn 186:16  c=7.17559e-17
c1363 364:cn 156:16  c=6.54455e-20
c1362 364:cn x27|src  c=4.20929e-20
c1361 364:cn 295:4  c=2.79154e-18
c1360 364:cn 187:16  c=1.77439e-17
c1359 364:cn m5|x1|drn  c=3.19267e-19
cg1358 363:cn gnd  c=2.34526e-17
c1357 363:cn 133:c  c=7.17966e-19
c1356 363:cn 137:14  c=5.48004e-18
c1355 363:cn 74:c  c=8.23915e-18
c1354 363:cn 82:c  c=8.83841e-17
c1353 363:cn 83:c  c=4.64693e-18
c1352 363:cn 32:rn  c=6.92865e-18
c1351 363:cn x2|src  c=6.23057e-19
c1350 363:cn 348:2  c=1.46165e-17
cg1349 362:cn gnd  c=1.90181e-17
c1348 362:cn 187:16  c=1.37342e-19
c1347 362:cn 82:c  c=6.77152e-17
c1346 362:cn 32:rn  c=5.62726e-18
c1345 362:cn 76:c  c=2.79504e-19
c1344 362:cn m18|x1|src  c=3.43005e-19
c1343 362:cn 118:c  c=5.35495e-18
c1342 362:cn 50:rn  c=4.66164e-19
c1341 362:cn 249:4  c=7.80593e-18
c1340 362:cn 285:4  c=8.2418e-19
c1339 362:cn 186:16  c=8.70544e-18
c1338 362:cn 156:16  c=1.09236e-18
cg1337 m11|x1|gate gnd  c=4.35279e-19
c1336 m11|x1|gate 338:2  c=1.36612e-18
c1335 m11|x1|gate 322:2  c=7.07278e-18
c1334 m11|x1|gate 216:9  c=9.0728e-20
c1333 m11|x1|gate 310:2  c=1.16212e-20
cg1332 359:cn gnd  c=3.4873e-18
c1331 359:cn 25:rn  c=4.84754e-21
c1330 359:cn x10|drn  c=5.59444e-19
c1329 359:cn x11|drn  c=5.68303e-19
c1328 359:cn 202:9  c=2.62301e-18
c1327 359:cn 293:4  c=3.82845e-18
c1326 359:cn 208:9  c=1.98324e-18
c1325 359:cn 269:4  c=1.98683e-18
cg1324 356:cn gnd  c=4.16669e-18
c1323 356:cn 216:9  c=2.07201e-18
c1322 356:cn x11|drn  c=5.68024e-19
c1321 356:cn x12|src  c=6.88178e-19
c1320 356:cn 293:4  c=4.10824e-18
c1319 356:cn 239:9  c=3.07065e-18
c1318 356:cn 322:2  c=6.88797e-22
c1317 356:cn 338:2  c=3.34507e-19
c1316 356:cn 84:c  c=1.51782e-20
c1315 356:cn 43:rn  c=4.79736e-21
c1314 356:cn 269:4  c=1.98709e-18
cg1313 355:cn gnd  c=1.69702e-17
c1312 355:cn 187:16  c=1.47499e-19
c1311 355:cn 250:4  c=2.99361e-18
c1310 355:cn 251:4  c=5.05583e-18
c1309 355:cn 82:c  c=8.83005e-17
c1308 355:cn 205:9  c=6.64991e-20
c1307 355:cn 32:rn  c=6.92865e-18
c1306 355:cn 81:c  c=3.73009e-18
c1305 355:cn 186:16  c=6.24588e-18
cg1304 354:cn gnd  c=8.09352e-17
c1303 354:cn 230:9  c=3.41857e-19
c1302 354:cn 203:9  c=3.61115e-19
c1301 354:cn 216:9  c=4.78777e-19
c1300 354:cn 6:rn  c=1.94212e-21
c1299 354:cn 232:9  c=9.00108e-20
c1298 354:cn 8:rn  c=2.58949e-21
c1297 354:cn 202:9  c=9.86793e-19
c1296 354:cn 250:4  c=2.25596e-19
c1295 354:cn 251:4  c=8.04233e-20
c1294 354:cn 239:9  c=4.43171e-19
c1293 354:cn 322:2  c=2.18986e-17
c1292 354:cn 205:9  c=6.1488e-18
c1291 354:cn 82:c  c=7.08611e-20
c1290 354:cn m11|x1|src  c=2.88117e-18
c1289 354:cn 131:c  c=1.08462e-17
c1288 354:cn 32:rn  c=7.08611e-20
c1287 354:cn 338:2  c=1.46171e-17
c1286 354:cn 310:2  c=1.76106e-17
c1285 354:cn 349:2  c=3.66932e-17
c1284 354:cn 51:rn  c=2.05733e-18
c1283 354:cn 84:c  c=8.72554e-18
c1282 354:cn 237:9  c=4.32984e-19
c1281 354:cn 86:c  c=1.1538e-17
c1280 354:cn 206:9  c=2.02571e-19
c1279 354:cn 77:c  c=3.18346e-20
c1278 354:cn 89:c  c=1.51673e-18
c1277 354:cn 40:rn  c=3.60054e-18
c1276 354:cn 27:rn  c=2.54927e-19
c1275 354:cn 43:rn  c=1.63258e-17
c1274 354:cn 44:rn  c=3.73234e-18
c1273 354:cn 45:rn  c=7.01779e-18
c1272 354:cn 41:rn  c=1.14526e-17
cg1271 353:2 gnd  c=3.43627e-18
c1270 353:2 198:9  c=1.53915e-19
c1269 353:2 232:9  c=4.63112e-21
c1268 353:2 32:rn  c=7.66906e-18
c1267 353:2 240:9  c=1.50441e-17
c1266 353:2 206:9  c=1.78971e-17
c1265 353:2 207:9  c=1.02181e-17
c1264 353:2 88:c  c=4.23174e-19
c1263 353:2 136:14  c=3.21944e-18
c1262 352:2 133:c  c=6.18374e-19
c1261 352:2 140:14  c=9.74846e-19
c1260 352:2 144:14  c=1.44535e-19
c1259 352:2 x26|src  c=8.601e-20
c1258 352:2 135:14  c=6.99179e-17
c1257 352:2 125:c  c=1.10309e-19
c1256 352:2 128:c  c=1.18027e-17
c1255 352:2 107:c  c=4.83812e-18
c1254 352:2 108:c  c=2.43564e-18
c1253 352:2 130:c  c=4.98839e-18
c1252 352:2 109:c  c=2.51362e-18
c1251 352:2 116:c  c=4.37079e-18
c1250 352:2 138:14  c=9.2409e-19
c1249 352:2 73:c  c=4.20191e-18
c1248 352:2 136:14  c=1.05979e-16
cg1247 351:2 gnd  c=8.18975e-18
c1246 351:2 220:9  c=1.98763e-18
c1245 351:2 x28|drn  c=5.67946e-19
c1244 351:2 125:c  c=1.0907e-18
c1243 351:2 240:9  c=3.50908e-18
cg1242 350:2 gnd  c=2.01678e-17
c1241 350:2 240:9  c=2.03712e-19
c1240 350:2 136:14  c=2.09018e-18
cg1239 349:2 gnd  c=1.3931e-17
c1238 349:2 46:rn  c=1.52182e-18
c1237 349:2 31:rn  c=2.39914e-18
c1236 349:2 39:rn  c=1.52182e-18
c1235 349:2 203:9  c=7.96584e-18
c1234 349:2 212:9  c=6.96976e-20
c1233 349:2 215:9  c=1.97452e-18
c1232 349:2 200:9  c=4.38365e-17
c1231 349:2 204:9  c=8.21853e-19
c1230 349:2 202:9  c=4.78184e-19
c1229 349:2 205:9  c=1.6508e-17
c1228 349:2 82:c  c=3.40064e-17
c1227 349:2 235:9  c=1.37008e-17
c1226 349:2 131:c  c=5.97414e-17
c1225 349:2 32:rn  c=3.56582e-17
c1224 349:2 51:rn  c=7.62625e-17
c1223 349:2 84:c  c=5.05797e-19
c1222 349:2 86:c  c=3.93257e-18
c1221 349:2 238:9  c=3.57214e-19
c1220 349:2 104:c  c=6.22268e-18
c1219 349:2 105:c  c=3.74612e-18
c1218 349:2 206:9  c=4.85606e-19
c1217 349:2 77:c  c=9.07311e-18
c1216 349:2 207:9  c=4.25768e-18
c1215 349:2 87:c  c=4.5486e-18
c1214 349:2 236:9  c=3.58979e-18
c1213 349:2 81:c  c=6.81534e-18
c1212 349:2 44:rn  c=8.35994e-19
c1211 349:2 45:rn  c=4.42394e-18
c1210 349:2 41:rn  c=3.49618e-17
c1209 349:2 m7|x1|drn  c=1.28786e-19
cg1208 348:2 gnd  c=6.24621e-17
c1207 348:2 133:c  c=2.98502e-17
c1206 348:2 140:14  c=8.70301e-20
c1205 348:2 137:14  c=5.23258e-17
c1204 348:2 x24|drn  c=1.13835e-19
c1203 348:2 74:c  c=6.37694e-18
c1202 348:2 82:c  c=3.65669e-17
c1201 348:2 142:14  c=9.27002e-19
c1200 348:2 x26|src  c=1.02125e-19
c1199 348:2 32:rn  c=3.70499e-18
c1198 348:2 135:14  c=1.32944e-19
c1197 348:2 128:c  c=6.87199e-20
c1196 348:2 207:9  c=3.07151e-17
c1195 348:2 x2|drn  c=5.71047e-19
c1194 348:2 88:c  c=2.84046e-19
c1193 348:2 126:c  c=4.62108e-18
c1192 348:2 136:14  c=1.03525e-17
cg1191 347:2 gnd  c=1.60137e-18
c1190 347:2 32:rn  c=1.09013e-18
c1189 347:2 125:c  c=6.14848e-18
c1188 347:2 106:c  c=2.51028e-18
c1187 347:2 240:9  c=2.64608e-18
c1186 347:2 128:c  c=4.10643e-18
c1185 347:2 107:c  c=1.17303e-19
c1184 347:2 138:14  c=9.65568e-19
c1183 347:2 136:14  c=5.46746e-17
c1182 346:2 221:9  c=1.7878e-17
c1181 346:2 234:9  c=3.1987e-20
c1180 346:2 207:9  c=2.36818e-18
cg1179 345:2 gnd  c=1.08516e-19
c1178 345:2 m5|x1|drn  c=4.18252e-20
c1177 345:2 207:9  c=1.07377e-19
c1176 345:2 221:9  c=3.26884e-19
c1175 345:2 234:9  c=1.45395e-21
cg1174 342:2 gnd  c=3.43256e-18
c1173 342:2 231:9  c=6.81959e-20
c1172 342:2 234:9  c=2.40996e-19
c1171 342:2 221:9  c=2.07466e-18
c1170 342:2 238:9  c=5.14232e-19
c1169 342:2 207:9  c=3.26893e-18
c1168 342:2 m5|x1|drn  c=6.98597e-19
cg1167 341:2 gnd  c=1.54966e-17
c1166 341:2 133:c  c=2.24455e-19
c1165 341:2 203:9  c=1.79745e-18
c1164 341:2 233:9  c=1.14852e-18
c1163 341:2 234:9  c=5.05256e-20
c1162 341:2 82:c  c=1.55641e-19
c1161 341:2 221:9  c=1.74897e-18
c1160 341:2 238:9  c=3.894e-19
c1159 341:2 207:9  c=4.48721e-17
c1158 341:2 m5|x1|drn  c=6.63033e-19
c1157 341:2 88:c  c=5.49055e-20
c1156 341:2 41:rn  c=2.2623e-20
c1155 341:2 126:c  c=2.56975e-19
cg1154 340:2 gnd  c=8.04871e-18
c1153 340:2 230:9  c=5.5013e-21
c1152 340:2 220:9  c=1.98763e-18
c1151 340:2 x28|drn  c=5.67946e-19
c1150 340:2 240:9  c=3.53734e-18
cg1149 339:2 gnd  c=8.19702e-18
c1148 339:2 218:9  c=2.05008e-18
c1147 339:2 230:9  c=6.66465e-19
c1146 339:2 198:9  c=3.87498e-18
c1145 339:2 x27|src  c=6.66715e-19
c1144 339:2 40:rn  c=5.5013e-21
cg1143 338:2 gnd  c=9.2579e-18
c1142 338:2 198:9  c=1.07907e-19
c1141 338:2 216:9  c=2.45103e-18
c1140 338:2 202:9  c=4.25052e-19
c1139 338:2 239:9  c=5.15319e-17
c1138 338:2 237:9  c=9.6613e-19
c1137 338:2 43:rn  c=1.27137e-19
cg1136 337:2 gnd  c=2.33796e-18
c1135 337:2 203:9  c=5.32272e-21
c1134 337:2 32:rn  c=6.82485e-18
c1133 337:2 51:rn  c=1.76074e-20
c1132 337:2 207:9  c=3.4286e-17
c1131 337:2 88:c  c=4.828e-20
c1130 336:2 198:9  c=2.36818e-18
c1129 336:2 218:9  c=1.77931e-17
cg1128 331:2 gnd  c=6.79291e-18
c1127 331:2 137:14  c=8.76575e-19
c1126 331:2 142:14  c=8.05107e-19
c1125 331:2 x2|drn  c=8.64146e-19
cg1124 329:2 gnd  c=5.87088e-18
c1123 329:2 140:14  c=8.05107e-19
c1122 329:2 x24|drn  c=8.62903e-19
c1121 329:2 x26|src  c=8.63311e-19
c1120 329:2 135:14  c=7.34475e-19
c1119 329:2 128:c  c=2.26778e-17
c1118 329:2 107:c  c=1.98621e-18
c1117 329:2 108:c  c=1.75643e-17
c1116 329:2 130:c  c=1.98778e-18
c1115 329:2 109:c  c=1.75605e-17
c1114 329:2 116:c  c=1.98778e-18
c1113 329:2 138:14  c=8.05107e-19
c1112 329:2 73:c  c=1.98621e-18
c1111 329:2 136:14  c=1.49393e-18
cg1110 328:2 gnd  c=4.95158e-18
c1109 328:2 220:9  c=1.98763e-18
c1108 328:2 x28|drn  c=5.67946e-19
c1107 328:2 128:c  c=7.0911e-19
c1106 328:2 240:9  c=3.16539e-18
c1105 327:2 240:9  c=2.34427e-18
c1104 327:2 220:9  c=1.75774e-17
c1103 326:2 240:9  c=2.36818e-18
c1102 326:2 220:9  c=1.75774e-17
cg1101 325:2 gnd  c=4.95334e-18
c1100 325:2 230:9  c=7.08489e-19
c1099 325:2 218:9  c=2.07323e-18
c1098 325:2 198:9  c=3.75683e-18
c1097 325:2 234:9  c=3.67992e-22
c1096 325:2 x27|src  c=6.97923e-19
c1095 325:2 43:rn  c=5.85327e-21
cg1094 322:2 gnd  c=8.64814e-18
c1093 322:2 216:9  c=6.35179e-18
c1092 322:2 239:9  c=2.93004e-18
c1091 322:2 86:c  c=2.33033e-19
cg1090 321:2 gnd  c=6.80602e-18
c1089 321:2 46:rn  c=1.04103e-18
c1088 321:2 39:rn  c=1.84868e-19
c1087 321:2 215:9  c=1.56789e-18
c1086 321:2 122:c  c=8.88116e-21
c1085 321:2 235:9  c=1.74484e-18
c1084 321:2 104:c  c=2.10374e-18
c1083 321:2 105:c  c=1.81243e-17
c1082 321:2 77:c  c=2.21409e-17
c1081 321:2 87:c  c=2.5063e-18
c1080 321:2 m7|x1|drn  c=5.39429e-19
c1079 321:2 41:rn  c=1.84868e-19
cg1078 319:2 gnd  c=3.31966e-17
c1077 319:2 144:14  c=2.33761e-19
c1076 319:2 74:c  c=4.65078e-18
c1075 319:2 82:c  c=1.01272e-18
c1074 319:2 32:rn  c=2.74001e-17
c1073 319:2 135:14  c=7.07062e-18
c1072 319:2 136:14  c=1.43797e-17
cg1071 312:2 gnd  c=9.02777e-18
c1070 312:2 x24|drn  c=8.63235e-19
c1069 312:2 125:c  c=2.05045e-18
c1068 312:2 106:c  c=1.77784e-17
c1067 312:2 128:c  c=2.05045e-18
c1066 312:2 138:14  c=8.05107e-19
c1065 312:2 136:14  c=7.48044e-19
cg1064 311:2 gnd  c=1.3661e-17
c1063 311:2 133:c  c=1.31269e-18
c1062 311:2 137:14  c=1.14999e-18
c1061 311:2 82:c  c=2.49566e-17
c1060 311:2 20:rn  c=6.13513e-20
c1059 311:2 32:rn  c=3.91714e-17
c1058 311:2 51:rn  c=2.52628e-20
c1057 311:2 135:14  c=4.17718e-19
c1056 311:2 128:c  c=4.8369e-18
c1055 311:2 240:9  c=9.49091e-19
c1054 311:2 206:9  c=8.00856e-19
c1053 311:2 207:9  c=5.17566e-17
c1052 311:2 88:c  c=4.93434e-18
c1051 311:2 136:14  c=5.89301e-17
c1050 310:2 230:9  c=2.81399e-19
c1049 310:2 198:9  c=9.2926e-20
c1048 310:2 232:9  c=5.11481e-19
c1047 310:2 202:9  c=2.22568e-17
c1046 310:2 239:9  c=1.05827e-17
c1045 310:2 205:9  c=8.88227e-18
c1044 310:2 131:c  c=2.04743e-18
c1043 310:2 32:rn  c=3.7997e-19
c1042 310:2 51:rn  c=5.6103e-18
c1041 310:2 84:c  c=6.81752e-20
c1040 310:2 237:9  c=3.72385e-18
c1039 310:2 86:c  c=1.75854e-19
c1038 310:2 12:rn  c=7.25327e-20
c1037 310:2 206:9  c=7.07555e-18
c1036 310:2 43:rn  c=5.52463e-18
c1035 310:2 81:c  c=1.85141e-19
c1034 310:2 44:rn  c=2.8558e-18
cg1033 308:2 gnd  c=1.00733e-17
c1032 308:2 203:9  c=4.69162e-19
c1031 308:2 232:9  c=6.31262e-20
c1030 308:2 206:9  c=1.91926e-18
c1029 308:2 207:9  c=1.43638e-17
c1028 308:2 44:rn  c=1.8295e-21
c1027 308:2 45:rn  c=7.17107e-21
c1026 308:2 88:c  c=4.98545e-19
c1025 x24|src 128:c  c=6.98359e-19
c1024 x24|src 125:c  c=6.98359e-19
c1023 x24|src 32:rn  c=5.70616e-20
c1022 x24|src 138:14  c=7.8002e-19
c1021 x24|src 136:14  c=1.19445e-19
c1020 x24|src 82:c  c=4.68765e-20
cg1019 307:2 gnd  c=2.04473e-17
c1018 307:2 144:14  c=5.72833e-19
c1017 307:2 82:c  c=7.62379e-18
c1016 307:2 x26|src  c=4.73309e-19
c1015 307:2 32:rn  c=4.46322e-17
c1014 307:2 135:14  c=4.92481e-18
c1013 307:2 240:9  c=8.34341e-19
c1012 307:2 136:14  c=2.83815e-17
cg1011 306:2 gnd  c=6.59902e-17
c1010 306:2 31:rn  c=6.91137e-18
c1009 306:2 198:9  c=1.96081e-17
c1008 306:2 239:9  c=2.13117e-18
c1007 306:2 82:c  c=6.94951e-18
c1006 306:2 32:rn  c=1.02523e-16
c1005 306:2 x27|src  c=3.81374e-19
c1004 306:2 x28|drn  c=4.35045e-19
c1003 306:2 237:9  c=3.96258e-18
c1002 306:2 12:rn  c=2.49065e-18
c1001 306:2 240:9  c=1.90977e-17
c1000 306:2 206:9  c=5.42543e-18
c999 306:2 207:9  c=1.95431e-18
c998 306:2 43:rn  c=4.42882e-20
c997 306:2 136:14  c=1.4406e-18
cg996 305:2 gnd  c=2.35862e-18
c995 305:2 31:rn  c=8.31827e-17
c994 305:2 198:9  c=2.26897e-18
c993 305:2 202:9  c=3.03942e-18
c992 305:2 239:9  c=3.1745e-18
c991 305:2 82:c  c=2.8093e-17
c990 305:2 32:rn  c=2.23824e-16
c989 305:2 51:rn  c=9.77654e-18
c988 305:2 237:9  c=7.80824e-18
c987 305:2 1:rn  c=1.21129e-19
c986 305:2 12:rn  c=4.47476e-18
c985 305:2 240:9  c=2.2558e-18
c984 305:2 206:9  c=5.53646e-17
c983 305:2 207:9  c=5.7071e-18
c982 305:2 43:rn  c=7.67662e-19
c981 305:2 44:rn  c=9.86994e-20
c980 305:2 136:14  c=7.87731e-19
cg979 304:2 gnd  c=7.42974e-18
c978 304:2 31:rn  c=1.22496e-17
c977 304:2 202:9  c=2.58472e-18
c976 304:2 82:c  c=9.30443e-19
c975 304:2 205:9  c=2.13002e-18
c974 304:2 32:rn  c=8.97649e-17
c973 304:2 1:rn  c=1.72976e-18
c972 304:2 12:rn  c=2.69495e-18
c971 304:2 206:9  c=5.50909e-20
c970 304:2 81:c  c=7.35629e-18
cg969 x2|src gnd  c=4.90839e-20
c968 x2|src 137:14  c=2.25602e-19
c967 x2|src 142:14  c=7.76216e-19
cg966 303:2 gnd  c=2.06449e-17
c965 303:2 230:9  c=7.59339e-19
c964 303:2 198:9  c=5.94899e-18
c963 303:2 234:9  c=8.40506e-21
c962 303:2 220:9  c=2.23922e-17
c961 303:2 221:9  c=8.57435e-20
c960 303:2 x28|drn  c=2.31608e-18
c959 303:2 238:9  c=1.26781e-19
c958 303:2 128:c  c=8.79518e-19
c957 303:2 240:9  c=1.75203e-17
c956 303:2 206:9  c=1.9451e-17
c955 303:2 m5|x1|drn  c=4.55705e-20
c954 303:2 43:rn  c=6.33547e-21
cg953 302:2 gnd  c=5.44776e-18
c952 302:2 230:9  c=8.41898e-23
c951 302:2 232:9  c=4.6917e-21
c950 302:2 240:9  c=1.1409e-19
c949 302:2 206:9  c=4.29412e-19
c948 302:2 207:9  c=8.87366e-20
c947 302:2 88:c  c=1.77361e-19
c946 302:2 136:14  c=4.9528e-19
cg945 300:2 gnd  c=7.33382e-18
c944 300:2 232:9  c=9.84685e-20
c943 300:2 206:9  c=4.31425e-18
c942 300:2 88:c  c=1.38063e-19
c941 300:2 136:14  c=4.4977e-19
c940 m7|x1|src 39:rn  c=1.0201e-19
c939 m7|x1|src 200:9  c=3.55895e-19
c938 m7|x1|src 204:9  c=1.17376e-19
c937 m7|x1|src 231:9  c=1.17376e-19
c936 m7|x1|src 104:c  c=4.29116e-19
c935 m7|x1|src 87:c  c=4.29116e-19
c934 m7|x1|src 77:c  c=2.65992e-18
c933 m7|x1|src 41:rn  c=1.0201e-19
cg932 297:2 gnd  c=5.00706e-18
c931 297:2 230:9  c=7.35327e-20
c930 297:2 198:9  c=2.75209e-19
c929 297:2 232:9  c=5.80759e-20
c928 297:2 237:9  c=3.69563e-20
c927 297:2 240:9  c=3.86652e-18
c926 297:2 206:9  c=1.57868e-18
c925 297:2 88:c  c=6.55808e-20
cg924 296:2 gnd  c=1.44373e-19
c923 296:2 230:9  c=5.85327e-21
c922 296:2 220:9  c=1.98763e-18
c921 296:2 x28|drn  c=5.67946e-19
c920 296:2 240:9  c=3.15233e-18
c919 x25|drn 133:c  c=9.07357e-20
c918 x25|drn 140:14  c=8.69213e-19
c917 x25|drn 74:c  c=3.87764e-20
c916 x25|drn 32:rn  c=1.35254e-20
c915 x25|drn 135:14  c=5.52344e-20
c914 x25|drn 128:c  c=3.05301e-18
c913 x25|drn 107:c  c=5.68958e-19
c912 x25|drn 130:c  c=5.67278e-19
c911 x25|drn 138:14  c=8.64665e-19
c910 x25|drn 116:c  c=5.67278e-19
c909 x25|drn 73:c  c=5.68958e-19
c908 x25|drn 136:14  c=9.44441e-20
c907 m11|x1|src 200:9  c=6.39843e-21
c906 m11|x1|src 131:c  c=8.14817e-20
c905 m11|x1|src 86:c  c=5.22003e-20
c904 m11|x1|src 81:c  c=3.14414e-20
cg903 295:4 gnd  c=6.73396e-18
c902 295:4 5:rn  c=3.74781e-18
c901 295:4 82:c  c=1.48099e-17
c900 295:4 32:rn  c=1.44416e-17
c899 295:4 155:16  c=6.37538e-19
c898 295:4 183:16  c=1.52943e-18
c897 295:4 157:16  c=1.19392e-18
c896 295:4 186:16  c=2.45851e-17
c895 295:4 156:16  c=5.74721e-18
cg894 294:4 gnd  c=2.32326e-17
c893 294:4 202:9  c=1.86239e-18
c892 293:4 216:9  c=9.52305e-19
c891 293:4 202:9  c=1.08e-16
c890 293:4 x12|src  c=1.01488e-19
c889 293:4 239:9  c=6.42241e-17
c888 293:4 208:9  c=9.43871e-19
cg887 292:4 gnd  c=6.92499e-18
c886 292:4 147:16  c=3.53734e-18
c885 292:4 33:rn  c=5.80175e-18
c884 292:4 23:rn  c=1.09856e-19
c883 292:4 x19|src  c=5.67946e-19
c882 292:4 169:16  c=1.98763e-18
cg881 291:4 gnd  c=9.55845e-19
c880 291:4 215:9  c=7.78453e-19
c879 291:4 187:16  c=3.36205e-18
c878 291:4 200:9  c=6.38528e-18
c877 291:4 158:16  c=6.81278e-19
c876 291:4 120:c  c=6.08642e-19
c875 291:4 205:9  c=3.00988e-19
c874 291:4 122:c  c=1.73568e-18
c873 291:4 235:9  c=2.69865e-17
c872 291:4 121:c  c=8.91218e-19
c871 291:4 236:9  c=6.65418e-19
cg870 290:4 gnd  c=6.59959e-18
c869 290:4 182:16  c=1.1985e-17
c868 290:4 146:16  c=3.09554e-18
c867 290:4 147:16  c=5.82695e-19
c866 290:4 118:c  c=1.51233e-18
c865 290:4 50:rn  c=6.16704e-18
c864 290:4 157:16  c=4.15956e-17
c863 290:4 103:c  c=1.87712e-18
c862 290:4 156:16  c=8.17529e-19
cg861 289:4 gnd  c=8.94865e-19
c860 289:4 25:rn  c=1.49493e-19
c859 289:4 202:9  c=5.03233e-17
c858 289:4 151:16  c=2.59297e-18
c857 289:4 208:9  c=9.3977e-19
c856 289:4 49:rn  c=7.6021e-19
c855 288:4 5:rn  c=2.78988e-17
c854 288:4 187:16  c=1.67957e-18
c853 288:4 158:16  c=8.05107e-19
c852 288:4 155:16  c=2.50182e-19
c851 288:4 185:16  c=2.01773e-21
c850 288:4 186:16  c=5.13666e-19
cg849 287:4 gnd  c=7.13629e-18
c848 287:4 4:rn  c=4.82033e-19
c847 287:4 5:rn  c=2.6463e-17
c846 287:4 146:16  c=1.12806e-19
c845 287:4 184:16  c=9.21926e-19
c844 287:4 183:16  c=3.05109e-18
c843 287:4 157:16  c=1.36953e-18
c842 287:4 186:16  c=2.71611e-18
c841 287:4 156:16  c=2.65551e-18
cg840 286:4 gnd  c=1.9836e-17
c839 286:4 5:rn  c=1.27012e-16
c838 286:4 187:16  c=1.5456e-18
c837 286:4 82:c  c=4.25167e-19
c836 286:4 155:16  c=8.92843e-18
c835 286:4 183:16  c=7.8019e-20
c834 286:4 186:16  c=2.89816e-17
c833 286:4 156:16  c=6.44771e-19
cg832 285:4 gnd  c=3.41126e-17
c831 285:4 182:16  c=1.63226e-18
c830 285:4 187:16  c=9.23633e-20
c829 285:4 146:16  c=7.54309e-18
c828 285:4 149:16  c=2.41219e-17
c827 285:4 82:c  c=4.71844e-18
c826 285:4 32:rn  c=4.01684e-18
c825 285:4 76:c  c=3.86964e-18
c824 285:4 153:16  c=5.99509e-18
c823 285:4 155:16  c=2.12911e-18
c822 285:4 118:c  c=2.76991e-17
c821 285:4 50:rn  c=3.61566e-17
c820 285:4 184:16  c=1.32624e-17
c819 285:4 183:16  c=9.78806e-19
c818 285:4 132:c  c=2.73946e-17
c817 285:4 75:c  c=7.62615e-19
c816 285:4 157:16  c=8.66629e-18
c815 285:4 103:c  c=1.42121e-18
c814 285:4 186:16  c=3.51536e-18
c813 285:4 156:16  c=3.64928e-18
c812 285:4 111:c  c=1.03056e-19
cg811 284:4 gnd  c=2.10003e-18
c810 284:4 37:rn  c=1.44818e-17
c809 284:4 187:16  c=7.2527e-19
c808 284:4 185:16  c=7.62562e-19
cg807 283:4 gnd  c=3.84301e-18
c806 283:4 4:rn  c=2.08577e-19
c805 283:4 5:rn  c=2.19026e-17
c804 283:4 48:rn  c=1.72829e-19
c803 283:4 8:rn  c=1.35484e-19
c802 283:4 146:16  c=3.16546e-19
c801 283:4 157:16  c=4.7343e-18
c800 283:4 156:16  c=1.00002e-18
cg799 281:4 gnd  c=2.31042e-17
c798 281:4 4:rn  c=5.45237e-18
c797 281:4 182:16  c=1.5923e-18
c796 281:4 146:16  c=3.2747e-18
c795 281:4 147:16  c=5.20851e-18
c794 281:4 151:16  c=2.68553e-19
c793 281:4 167:16  c=2.40298e-17
c792 281:4 x17|drn  c=3.13657e-18
c791 281:4 157:16  c=2.89962e-17
c790 281:4 103:c  c=3.0069e-22
cg789 279:4 gnd  c=5.20347e-18
c788 279:4 103:c  c=1.43825e-19
c787 279:4 157:16  c=2.59909e-18
c786 279:4 182:16  c=3.73428e-18
cg785 278:4 gnd  c=8.18119e-18
c784 278:4 167:16  c=1.98763e-18
c783 278:4 x17|drn  c=5.67946e-19
c782 278:4 165:16  c=2.63716e-20
c781 278:4 157:16  c=3.53734e-18
c780 278:4 188:16  c=6.66184e-19
cg779 277:4 gnd  c=1.45502e-17
c778 277:4 118:c  c=6.19034e-18
cg777 276:4 gnd  c=3.5018e-18
c776 276:4 3:rn  c=5.84213e-20
c775 276:4 22:rn  c=3.13813e-18
c774 276:4 147:16  c=2.70735e-18
c773 276:4 x19|src  c=5.67946e-19
c772 276:4 169:16  c=1.98763e-18
cg771 270:4 gnd  c=1.44955e-17
c770 270:4 x1|src  c=8.79945e-19
c769 270:4 215:9  c=8.05107e-19
c768 270:4 5:rn  c=1.2569e-19
c767 270:4 37:rn  c=4.50026e-19
c766 270:4 187:16  c=5.35843e-18
c765 270:4 200:9  c=1.61745e-18
c764 270:4 158:16  c=5.3016e-19
c763 270:4 120:c  c=2.07345e-18
c762 270:4 122:c  c=1.83591e-17
c761 270:4 235:9  c=1.66617e-17
c760 270:4 121:c  c=4.12962e-18
c759 270:4 77:c  c=1.97929e-19
c758 270:4 87:c  c=6.6937e-19
cg757 269:4 gnd  c=6.67556e-18
c756 269:4 x10|drn  c=8.6306e-19
c755 269:4 216:9  c=8.05107e-19
c754 269:4 202:9  c=1.4601e-18
c753 269:4 x12|src  c=7.75302e-19
c752 269:4 239:9  c=7.69922e-19
c751 269:4 208:9  c=8.05107e-19
c750 268:4 34:rn  c=5.09855e-19
c749 268:4 147:16  c=2.36818e-18
c748 268:4 169:16  c=1.75774e-17
c747 267:4 167:16  c=1.75774e-17
c746 267:4 157:16  c=2.36818e-18
cg745 266:4 gnd  c=8.04871e-18
c744 266:4 167:16  c=1.98763e-18
c743 266:4 x17|drn  c=5.67946e-19
c742 266:4 33:rn  c=1.09856e-19
c741 266:4 157:16  c=3.53734e-18
c740 266:4 188:16  c=5.5013e-21
cg739 264:4 gnd  c=6.52677e-18
c738 264:4 146:16  c=6.32656e-21
c737 264:4 m18|x1|drn  c=5.39429e-19
c736 264:4 155:16  c=7.31294e-19
c735 264:4 185:16  c=7.38131e-20
c734 264:4 184:16  c=1.66777e-19
c733 263:4 167:16  c=1.75774e-17
c732 263:4 157:16  c=2.36818e-18
cg731 261:4 gnd  c=8.7793e-18
c730 261:4 181:16  c=6.57481e-19
c729 261:4 182:16  c=7.38131e-20
c728 261:4 145:16  c=1.52588e-21
c727 261:4 x9|drn  c=5.39429e-19
c726 261:4 153:16  c=1.73835e-19
c725 261:4 165:16  c=2.95389e-19
c724 261:4 166:16  c=1.82982e-19
c723 261:4 119:c  c=2.10197e-18
c722 261:4 102:c  c=1.80192e-17
c721 261:4 103:c  c=2.07332e-18
c720 261:4 188:16  c=7.38131e-20
cg719 259:4 gnd  c=4.00091e-17
c718 259:4 202:9  c=1.43713e-17
c717 259:4 239:9  c=5.75817e-18
c716 259:4 82:c  c=4.67576e-18
c715 259:4 32:rn  c=2.76419e-17
cg714 252:4 gnd  c=1.28164e-17
c713 252:4 25:rn  c=2.73439e-20
c712 252:4 x10|drn  c=8.63027e-19
c711 252:4 202:9  c=7.93763e-19
c710 252:4 208:9  c=8.05107e-19
c709 252:4 49:rn  c=2.73439e-20
c708 252:4 26:rn  c=2.43562e-19
cg707 251:4 gnd  c=1.01302e-18
c706 251:4 4:rn  c=7.62212e-19
c705 251:4 5:rn  c=6.19666e-18
c704 251:4 187:16  c=5.475e-18
c703 251:4 48:rn  c=9.07967e-17
c702 251:4 6:rn  c=3.52802e-18
c701 251:4 8:rn  c=5.63844e-18
c700 251:4 202:9  c=1.75733e-16
c699 251:4 146:16  c=2.7224e-19
c698 251:4 158:16  c=1.89035e-19
c697 251:4 120:c  c=2.23643e-18
c696 251:4 205:9  c=1.29516e-16
c695 251:4 82:c  c=3.17999e-17
c694 251:4 235:9  c=1.24659e-17
c693 251:4 131:c  c=2.57143e-18
c692 251:4 151:16  c=1.5494e-18
c691 251:4 32:rn  c=1.92878e-17
c690 251:4 123:c  c=6.51745e-19
c689 251:4 84:c  c=4.80626e-18
c688 251:4 86:c  c=2.66423e-19
c687 251:4 1:rn  c=4.5976e-18
c686 251:4 12:rn  c=1.33241e-18
c685 251:4 89:c  c=2.45697e-17
c684 251:4 157:16  c=8.06138e-17
c683 251:4 236:9  c=4.11256e-18
c682 251:4 186:16  c=1.27248e-18
c681 251:4 156:16  c=1.84145e-18
cg680 250:4 gnd  c=1.89044e-18
c679 250:4 5:rn  c=1.65285e-17
c678 250:4 187:16  c=7.51924e-19
c677 250:4 x5|drn  c=4.0917e-19
c676 250:4 48:rn  c=1.66664e-18
c675 250:4 202:9  c=6.26319e-18
c674 250:4 146:16  c=2.20939e-19
c673 250:4 158:16  c=2.59303e-19
c672 250:4 205:9  c=2.21749e-17
c671 250:4 82:c  c=4.05974e-17
c670 250:4 151:16  c=8.85259e-20
c669 250:4 32:rn  c=8.5921e-17
c668 250:4 84:c  c=2.73688e-19
c667 250:4 184:16  c=5.81304e-19
c666 250:4 183:16  c=1.34385e-18
c665 250:4 1:rn  c=5.16102e-18
c664 250:4 157:16  c=3.58293e-17
c663 250:4 186:16  c=2.14018e-17
c662 250:4 156:16  c=1.16857e-17
cg661 249:4 gnd  c=1.1826e-16
c660 249:4 155:16  c=2.00136e-18
c659 249:4 185:16  c=8.63332e-19
c658 249:4 184:16  c=4.93741e-18
c657 249:4 145:16  c=3.71362e-19
c656 249:4 146:16  c=1.09012e-18
c655 249:4 149:16  c=2.48357e-18
c654 249:4 x9|drn  c=1.98542e-19
c653 249:4 152:16  c=1.71874e-18
c652 249:4 75:c  c=6.71926e-18
c651 249:4 153:16  c=5.18595e-17
c650 249:4 154:16  c=1.9036e-18
c649 249:4 165:16  c=6.08357e-19
c648 249:4 119:c  c=4.60126e-18
c647 249:4 102:c  c=3.60849e-18
c646 249:4 103:c  c=4.68476e-17
c645 249:4 111:c  c=1.26128e-18
c644 249:4 188:16  c=8.15666e-19
c643 249:4 132:c  c=1.03263e-16
c642 249:4 181:16  c=8.15666e-19
c641 249:4 182:16  c=7.40457e-18
c640 249:4 157:16  c=5.79083e-18
c639 249:4 m18|x1|drn  c=1.68959e-19
c638 249:4 76:c  c=7.60584e-18
c637 249:4 118:c  c=3.21826e-17
c636 249:4 50:rn  c=5.86158e-17
c635 x10|src 208:9  c=7.77944e-19
c634 x10|src 202:9  c=1.21154e-19
c633 x9|src 188:16  c=1.85005e-19
c632 x9|src 119:c  c=4.03631e-19
c631 x9|src 182:16  c=1.85005e-19
c630 x9|src 103:c  c=3.74528e-19
c629 x9|src 153:16  c=9.02118e-20
cg628 247:4 gnd  c=3.6656e-17
c627 247:4 4:rn  c=7.7973e-17
c626 247:4 182:16  c=3.28545e-18
c625 247:4 5:rn  c=2.50237e-18
c624 247:4 48:rn  c=5.79537e-19
c623 247:4 6:rn  c=9.45073e-18
c622 247:4 8:rn  c=8.33745e-20
c621 247:4 171:16  c=4.80739e-19
c620 247:4 3:rn  c=2.08577e-19
c619 247:4 22:rn  c=2.08577e-19
c618 247:4 146:16  c=1.6674e-16
c617 247:4 147:16  c=4.93624e-18
c616 247:4 151:16  c=1.3191e-18
c615 247:4 167:16  c=7.14629e-19
c614 247:4 m18|x1|drn  c=2.37944e-20
c613 247:4 184:16  c=9.55273e-18
c612 247:4 183:16  c=1.62227e-19
c611 247:4 157:16  c=5.50369e-17
c610 247:4 169:16  c=6.09452e-18
c609 247:4 103:c  c=1.24649e-19
c608 247:4 186:16  c=1.29136e-18
c607 247:4 156:16  c=3.47339e-18
cg606 246:4 gnd  c=3.20811e-17
c605 246:4 48:rn  c=6.73114e-19
c604 246:4 202:9  c=2.75123e-17
c603 246:4 x12|src  c=1.33454e-19
c602 246:4 239:9  c=5.30795e-18
c601 246:4 82:c  c=6.39397e-18
c600 246:4 151:16  c=1.45037e-18
c599 246:4 32:rn  c=4.2292e-17
c598 246:4 12:rn  c=2.21671e-17
c597 m18|x1|src 155:16  c=1.85005e-19
c596 m18|x1|src 185:16  c=1.85005e-19
c595 m18|x1|src 184:16  c=2.99468e-19
c594 m18|x1|src 157:16  c=9.83853e-20
c593 x1|drn 236:9  c=1.35206e-19
c592 x1|drn 235:9  c=1.17546e-19
c591 x1|drn 121:c  c=7.25723e-19
c590 x1|drn 120:c  c=7.22467e-19
c589 x1|drn 215:9  c=7.75325e-19
c588 x1|drn 200:9  c=5.4068e-19
cg587 245:4 gnd  c=3.5018e-18
c586 245:4 182:16  c=4.79736e-21
c585 245:4 22:rn  c=5.84213e-20
c584 245:4 167:16  c=1.98763e-18
c583 245:4 x17|drn  c=5.67946e-19
c582 245:4 157:16  c=2.70735e-18
cg581 243:4 gnd  c=4.36488e-18
c580 243:4 182:16  c=1.95866e-20
c579 243:4 6:rn  c=3.89908e-20
c578 243:4 48:rn  c=8.31453e-21
c577 243:4 146:16  c=2.08577e-19
c576 243:4 2:rn  c=2.1529e-19
c575 243:4 147:16  c=2.29618e-18
c574 243:4 151:16  c=3.50488e-19
c573 243:4 157:16  c=1.0003e-17
c572 x11|drn 216:9  c=8.67193e-19
c571 x11|drn 202:9  c=1.38312e-19
c570 x11|drn 239:9  c=4.60327e-20
c569 x11|drn 208:9  c=8.66437e-19
c568 242:4 25:rn  c=2.04402e-19
c567 242:4 4:rn  c=5.93516e-19
c566 242:4 5:rn  c=4.53693e-19
c565 242:4 48:rn  c=7.56674e-17
c564 242:4 6:rn  c=2.04881e-18
c563 242:4 8:rn  c=2.64946e-18
c562 242:4 202:9  c=5.58053e-17
c561 242:4 2:rn  c=1.58887e-19
c560 242:4 239:9  c=5.42717e-19
c559 242:4 205:9  c=8.7767e-20
c558 242:4 151:16  c=5.81387e-19
c557 242:4 32:rn  c=2.11765e-18
c556 242:4 1:rn  c=1.39347e-18
c555 242:4 12:rn  c=9.93283e-18
c554 242:4 157:16  c=6.84401e-19
c553 242:4 156:16  c=3.27038e-21
c552 241:4 155:16  c=3.51825e-19
c551 241:4 118:c  c=5.59815e-19
c550 241:4 184:16  c=4.73259e-19
cg549 240:9 gnd  c=5.67462e-18
cg548 239:9 gnd  c=6.75513e-18
cg547 238:9 gnd  c=1.17058e-17
c546 238:9 82:c  c=4.2438e-18
c545 238:9 41:rn  c=1.05425e-19
cg544 237:9 gnd  c=5.98206e-18
c543 237:9 43:rn  c=4.30103e-18
cg542 236:9 gnd  c=8.06166e-18
c541 236:9 81:c  c=9.65301e-19
c540 236:9 82:c  c=3.74133e-18
cg539 235:9 gnd  c=1.24247e-18
c538 235:9 120:c  c=2.4592e-18
c537 235:9 122:c  c=2.47991e-18
c536 235:9 131:c  c=9.82245e-20
c535 235:9 121:c  c=4.87042e-18
c534 235:9 123:c  c=3.48731e-19
c533 235:9 84:c  c=8.57506e-19
c532 235:9 104:c  c=7.24594e-20
c531 235:9 87:c  c=3.68474e-19
c530 235:9 77:c  c=1.30993e-17
c529 235:9 89:c  c=1.275e-18
cg528 234:9 gnd  c=8.65517e-18
c527 234:9 39:rn  c=9.20639e-21
cg526 233:9 gnd  c=4.34594e-18
c525 233:9 41:rn  c=2.17407e-19
cg524 232:9 gnd  c=6.59271e-18
c523 232:9 51:rn  c=4.48645e-19
c522 232:9 43:rn  c=9.92894e-18
c521 232:9 44:rn  c=1.75994e-17
cg520 231:9 gnd  c=3.77974e-18
c519 231:9 39:rn  c=1.43613e-17
c518 231:9 87:c  c=4.77527e-19
cg517 230:9 gnd  c=2.02125e-17
c516 230:9 40:rn  c=3.57915e-18
c515 230:9 27:rn  c=5.09855e-19
c514 230:9 43:rn  c=1.46934e-17
c513 x1|src 120:c  c=7.27395e-19
c512 x1|src 121:c  c=7.27395e-19
c511 x1|src 123:c  c=3.76652e-21
c510 x1|src 84:c  c=5.14777e-19
c509 x1|src 77:c  c=2.60351e-18
cg508 221:9 gnd  c=6.57394e-18
cg507 220:9 gnd  c=5.47311e-18
cg506 218:9 gnd  c=8.18224e-18
cg505 216:9 gnd  c=1.27277e-17
c504 216:9 84:c  c=3.75337e-19
cg503 215:9 gnd  c=8.6888e-18
c502 215:9 120:c  c=2.07472e-18
c501 215:9 122:c  c=1.78652e-17
c500 215:9 121:c  c=2.07472e-18
c499 215:9 84:c  c=9.66026e-19
c498 215:9 105:c  c=2.71652e-20
c497 215:9 77:c  c=2.20765e-17
c496 215:9 87:c  c=4.02554e-19
cg495 212:9 gnd  c=2.84892e-17
c494 212:9 82:c  c=7.27483e-18
cg493 208:9 gnd  c=6.68213e-18
cg492 207:9 gnd  c=2.54145e-17
c491 207:9 31:rn  c=2.26888e-19
c490 207:9 82:c  c=3.669e-17
c489 207:9 131:c  c=9.91907e-21
c488 207:9 32:rn  c=3.11583e-17
c487 207:9 51:rn  c=1.15938e-18
c486 207:9 45:rn  c=1.22289e-19
cg485 206:9 gnd  c=1.54154e-17
c484 206:9 31:rn  c=3.9641e-18
c483 206:9 82:c  c=1.61732e-17
c482 206:9 32:rn  c=5.40828e-17
c481 206:9 51:rn  c=3.90528e-17
c480 206:9 43:rn  c=1.99019e-18
c479 206:9 44:rn  c=4.60951e-18
c478 206:9 45:rn  c=4.35111e-19
cg477 205:9 gnd  c=4.48024e-18
c476 205:9 48:rn  c=1.4714e-20
c475 205:9 120:c  c=5.92353e-19
c474 205:9 82:c  c=2.03791e-17
c473 205:9 131:c  c=8.34979e-17
c472 205:9 32:rn  c=3.45725e-17
c471 205:9 123:c  c=3.21457e-19
c470 205:9 51:rn  c=2.35474e-19
c469 205:9 84:c  c=2.0267e-17
c468 205:9 86:c  c=2.98165e-18
c467 205:9 12:rn  c=8.09585e-20
c466 205:9 104:c  c=1.48863e-19
c465 205:9 89:c  c=2.30591e-17
c464 205:9 81:c  c=4.72585e-18
c463 205:9 41:rn  c=1.92358e-19
cg462 204:9 gnd  c=5.93991e-18
c461 204:9 46:rn  c=1.39252e-17
c460 204:9 104:c  c=4.77527e-19
c459 204:9 105:c  c=4.77527e-19
c458 204:9 89:c  c=5.29697e-21
c457 204:9 41:rn  c=3.05567e-17
cg456 203:9 gnd  c=5.44693e-17
c455 203:9 82:c  c=4.25167e-19
c454 203:9 32:rn  c=4.25167e-19
c453 203:9 51:rn  c=1.17581e-17
c452 203:9 89:c  c=4.50806e-21
c451 203:9 44:rn  c=8.41527e-18
c450 203:9 45:rn  c=2.69978e-17
c449 203:9 41:rn  c=1.21297e-16
cg448 202:9 gnd  c=4.45084e-18
c447 202:9 48:rn  c=2.618e-18
c446 202:9 82:c  c=4.44325e-19
c445 202:9 32:rn  c=1.9759e-17
c444 202:9 84:c  c=1.60332e-18
c443 202:9 12:rn  c=1.95473e-18
cg442 200:9 gnd  c=5.21116e-17
c441 200:9 46:rn  c=3.34059e-19
c440 200:9 39:rn  c=1.74622e-19
c439 200:9 x6|src  c=6.79105e-19
c438 200:9 82:c  c=1.75223e-17
c437 200:9 104:c  c=3.79613e-21
c436 200:9 105:c  c=1.6703e-19
c435 200:9 87:c  c=8.7311e-20
c434 200:9 41:rn  c=1.47212e-21
c433 200:9 m7|x1|drn  c=6.79105e-19
c432 x27|src 82:c  c=2.03393e-20
c431 m10|x1|gate 27:rn  c=2.54927e-19
c430 x28|drn 82:c  c=1.31041e-20
c429 x28|drn 32:rn  c=7.41538e-20
cg428 198:9 gnd  c=8.36016e-18
c427 198:9 43:rn  c=8.2739e-20
cg426 196:q gnd  c=6.70949e-18
c425 196:q 145:16  c=1.98763e-18
c424 196:q 148:16  c=1.98763e-18
c423 196:q 152:16  c=2.25813e-17
c422 196:q 153:16  c=1.01429e-20
c421 196:q 163:16  c=1.98763e-18
c420 196:q 164:16  c=1.75774e-17
c419 196:q 165:16  c=1.98763e-18
c418 196:q 166:16  c=1.75774e-17
cg417 193:q gnd  c=7.74901e-18
c416 193:q 154:16  c=2.08225e-18
c415 193:q 161:16  c=1.7878e-17
c414 193:q 162:16  c=2.07466e-18
cg413 192:q gnd  c=1.53776e-17
c412 192:q 159:16  c=2.07466e-18
c411 192:q 160:16  c=1.7878e-17
c410 192:q 152:16  c=2.07466e-18
cg409 191:q gnd  c=1.27487e-16
c408 191:q 153:16  c=5.1702e-17
c407 191:q 154:16  c=2.10647e-17
c406 191:q 161:16  c=2.36818e-18
c405 191:q 162:16  c=3.29311e-18
c404 m23|x1|drn 162:16  c=7.43977e-19
c403 m23|x1|drn 154:16  c=7.40118e-19
c402 x13|src 159:16  c=7.43977e-19
c401 x13|src 152:16  c=7.43977e-19
cg400 190:q gnd  c=2.61821e-17
c399 190:q 145:16  c=2.70735e-18
c398 190:q 148:16  c=2.70735e-18
c397 190:q 152:16  c=2.09233e-17
c396 190:q 153:16  c=1.40862e-18
c395 190:q 163:16  c=3.53734e-18
c394 190:q 164:16  c=2.36818e-18
c393 190:q 165:16  c=3.53734e-18
c392 190:q 166:16  c=2.36818e-18
c391 x14|drn 145:16  c=5.67946e-19
c390 x14|drn 148:16  c=5.67946e-19
c389 x14|drn 152:16  c=2.64205e-18
c388 x14|drn 163:16  c=5.67946e-19
c387 x14|drn 165:16  c=5.67946e-19
cg386 189:q gnd  c=7.06611e-17
c385 189:q 159:16  c=3.96418e-18
c384 189:q 160:16  c=2.36818e-18
c383 189:q 152:16  c=2.84767e-17
c382 189:q 153:16  c=3.87623e-17
cg381 188:16 gnd  c=4.69175e-18
c380 188:16 119:c  c=1.43017e-17
cg379 187:16 gnd  c=1.1959e-17
c378 187:16 x4|src  c=2.96099e-19
c377 187:16 5:rn  c=2.24414e-17
c376 187:16 37:rn  c=2.60924e-18
cg375 186:16 gnd  c=2.42891e-17
c374 186:16 x4|src  c=6.09521e-19
c373 186:16 5:rn  c=2.02536e-17
c372 186:16 82:c  c=6.387e-17
c371 186:16 32:rn  c=1.12338e-17
c370 186:16 m18|x1|drn  c=1.75669e-19
c369 186:16 118:c  c=2.34595e-18
c368 186:16 50:rn  c=6.76126e-19
c367 186:16 132:c  c=6.07244e-20
cg366 185:16 gnd  c=1.92978e-18
c365 185:16 37:rn  c=1.17653e-20
cg364 184:16 gnd  c=1.60577e-17
c363 184:16 5:rn  c=9.2576e-21
c362 184:16 32:rn  c=9.02635e-20
c361 184:16 50:rn  c=3.28374e-19
c360 184:16 132:c  c=6.87163e-18
c359 184:16 75:c  c=3.98268e-18
c358 184:16 103:c  c=5.98843e-18
c357 184:16 111:c  c=9.95719e-20
cg356 183:16 gnd  c=3.36973e-18
c355 183:16 5:rn  c=3.39445e-20
cg354 182:16 gnd  c=9.41921e-18
c353 182:16 103:c  c=8.0286e-17
c352 181:16 102:c  c=1.38786e-17
c351 x5|drn 48:rn  c=1.24809e-19
c350 x5|drn 32:rn  c=1.18403e-19
c349 x5|drn 8:rn  c=1.39567e-19
cg348 171:16 gnd  c=7.35652e-18
c347 171:16 25:rn  c=1.98763e-18
c346 171:16 4:rn  c=2.22944e-17
c345 171:16 3:rn  c=1.98763e-18
c344 171:16 23:rn  c=1.98763e-18
c343 171:16 24:rn  c=1.75774e-17
c342 171:16 49:rn  c=1.98763e-18
c341 171:16 26:rn  c=1.75774e-17
cg340 169:16 gnd  c=8.51683e-18
c339 169:16 22:rn  c=1.98763e-18
c338 169:16 33:rn  c=1.98763e-18
c337 169:16 34:rn  c=1.75774e-17
cg336 167:16 gnd  c=6.70949e-18
cg335 165:16 gnd  c=8.18119e-18
c334 165:16 119:c  c=6.66184e-19
cg333 163:16 gnd  c=8.05661e-18
cg332 162:16 gnd  c=2.70741e-18
cg331 159:16 gnd  c=8.76437e-18
cg330 158:16 gnd  c=7.6311e-18
c329 158:16 x4|src  c=5.57673e-19
c328 158:16 5:rn  c=2.23245e-17
c327 158:16 6:rn  c=1.04401e-19
c326 158:16 8:rn  c=1.24951e-19
c325 158:16 120:c  c=8.31679e-20
cg324 157:16 gnd  c=1.6961e-17
c323 157:16 1:rn  c=1.62166e-18
c322 157:16 12:rn  c=6.54125e-18
c321 157:16 x4|src  c=5.99688e-21
c320 157:16 4:rn  c=1.23844e-17
c319 157:16 5:rn  c=2.41271e-18
c318 157:16 6:rn  c=2.72045e-18
c317 157:16 8:rn  c=3.89482e-19
c316 157:16 82:c  c=5.27052e-18
c315 157:16 32:rn  c=4.67548e-17
c314 157:16 2:rn  c=8.39598e-19
c313 157:16 118:c  c=5.57663e-18
c312 157:16 50:rn  c=2.89662e-17
c311 157:16 48:rn  c=2.63586e-17
cg310 156:16 gnd  c=4.66765e-18
c309 156:16 5:rn  c=8.55389e-20
c308 156:16 48:rn  c=5.7104e-20
c307 156:16 82:c  c=2.6826e-18
c306 156:16 32:rn  c=3.24119e-17
c305 156:16 50:rn  c=3.57037e-18
c304 156:16 1:rn  c=3.00251e-19
c303 156:16 12:rn  c=1.27434e-19
cg302 155:16 gnd  c=1.28363e-17
c301 155:16 5:rn  c=2.4041e-19
c300 155:16 75:c  c=4.12371e-21
cg299 154:16 gnd  c=9.565e-18
cg298 153:16 gnd  c=7.74899e-17
c297 153:16 132:c  c=1.11622e-17
c296 153:16 75:c  c=6.44061e-18
c295 153:16 103:c  c=9.26645e-19
c294 153:16 111:c  c=1.67744e-17
cg293 152:16 gnd  c=2.9317e-17
c292 152:16 103:c  c=1.04173e-18
cg291 151:16 gnd  c=8.73486e-18
c290 151:16 25:rn  c=2.71681e-18
c289 151:16 4:rn  c=1.70522e-17
c288 151:16 48:rn  c=1.82698e-17
c287 151:16 8:rn  c=2.41069e-19
c286 151:16 3:rn  c=2.70735e-18
c285 151:16 2:rn  c=3.48393e-18
c284 151:16 12:rn  c=4.75955e-18
c283 151:16 23:rn  c=3.53734e-18
c282 151:16 24:rn  c=2.36818e-18
c281 151:16 49:rn  c=3.50536e-18
c280 151:16 26:rn  c=2.34392e-18
cg279 149:16 gnd  c=8.20697e-18
c278 149:16 118:c  c=4.25167e-19
c277 149:16 50:rn  c=3.94798e-19
c276 149:16 132:c  c=1.16166e-17
c275 149:16 75:c  c=1.82832e-17
c274 149:16 103:c  c=1.02541e-17
c273 149:16 111:c  c=2.46126e-18
cg272 148:16 gnd  c=3.5018e-18
cg271 147:16 gnd  c=7.16745e-18
c270 147:16 4:rn  c=5.49464e-18
c269 147:16 48:rn  c=5.95434e-19
c268 147:16 22:rn  c=2.70735e-18
c267 147:16 2:rn  c=3.02711e-19
c266 147:16 33:rn  c=3.53734e-18
c265 147:16 34:rn  c=2.36818e-18
c264 147:16 12:rn  c=8.2382e-19
cg263 146:16 gnd  c=1.26096e-17
c262 146:16 5:rn  c=6.77463e-21
c261 146:16 75:c  c=1.79608e-19
c260 146:16 103:c  c=5.98847e-18
c259 x21|src 25:rn  c=5.67946e-19
c258 x21|src 4:rn  c=2.76211e-18
c257 x21|src 3:rn  c=5.67946e-19
c256 x21|src 23:rn  c=5.67946e-19
c255 x21|src 49:rn  c=5.67946e-19
c254 x19|src 22:rn  c=5.67946e-19
c253 x19|src 33:rn  c=5.67946e-19
cg252 145:16 gnd  c=4.18454e-18
c251 145:16 103:c  c=5.82173e-19
cg250 144:14 gnd  c=9.69746e-18
c249 144:14 61:d  c=3.51403e-18
c248 144:14 62:d  c=2.34815e-18
c247 144:14 72:d  c=1.25538e-17
c246 144:14 71:d  c=3.53734e-18
c245 144:14 63:d  c=2.36818e-18
c244 144:14 64:d  c=3.004e-18
c243 144:14 56:d  c=1.82706e-17
c242 144:14 58:d  c=2.50257e-18
c241 144:14 59:d  c=3.02578e-19
c240 144:14 53:d  c=3.01948e-18
c239 144:14 128:c  c=1.45744e-19
c238 144:14 54:d  c=4.01484e-18
c237 144:14 88:c  c=4.06192e-19
cg236 143:14 gnd  c=5.60422e-18
c235 143:14 61:d  c=1.98763e-18
c234 143:14 62:d  c=1.75774e-17
c233 143:14 71:d  c=1.98763e-18
c232 143:14 63:d  c=1.75774e-17
c231 143:14 64:d  c=1.98763e-18
c230 143:14 56:d  c=2.24088e-17
c229 143:14 53:d  c=1.98763e-18
cg228 142:14 gnd  c=7.10942e-18
c227 142:14 56:d  c=8.38437e-20
c226 142:14 57:d  c=1.9565e-17
c225 142:14 69:d  c=1.98763e-18
cg224 140:14 gnd  c=6.3404e-18
c223 140:14 66:d  c=1.75774e-17
c222 140:14 60:d  c=1.98763e-18
c221 140:14 130:c  c=1.98022e-18
c220 140:14 109:c  c=1.75407e-17
c219 140:14 116:c  c=1.98022e-18
c218 140:14 65:d  c=1.98763e-18
cg217 138:14 gnd  c=5.98387e-18
c216 138:14 125:c  c=1.98181e-18
c215 138:14 106:c  c=1.75473e-17
c214 138:14 128:c  c=2.44962e-17
c213 138:14 107:c  c=1.98425e-18
c212 138:14 108:c  c=1.75606e-17
c211 138:14 73:c  c=1.98425e-18
cg210 137:14 gnd  c=1.84397e-17
c209 137:14 133:c  c=6.81048e-18
c208 137:14 72:d  c=2.11161e-19
c207 137:14 134:c  c=1.77028e-17
c206 137:14 52:rn  c=1.52502e-17
c205 137:14 74:c  c=1.70004e-18
c204 137:14 82:c  c=3.52169e-17
c203 137:14 57:d  c=6.5379e-17
c202 137:14 69:d  c=2.9983e-18
c201 137:14 83:c  c=3.31183e-18
c200 137:14 20:rn  c=4.18393e-18
c199 137:14 32:rn  c=4.78867e-17
c198 137:14 88:c  c=4.96568e-18
c197 137:14 126:c  c=1.78543e-18
cg196 136:14 gnd  c=3.63602e-18
c195 136:14 133:c  c=2.8438e-17
c194 136:14 72:d  c=1.01544e-17
c193 136:14 52:rn  c=1.14025e-18
c192 136:14 74:c  c=3.1029e-18
c191 136:14 56:d  c=1.88461e-17
c190 136:14 82:c  c=1.26504e-17
c189 136:14 57:d  c=6.56996e-18
c188 136:14 20:rn  c=3.81427e-19
c187 136:14 32:rn  c=9.27236e-17
c186 136:14 58:d  c=4.48237e-18
c185 136:14 59:d  c=3.234e-19
c184 136:14 125:c  c=3.3337e-18
c183 136:14 106:c  c=2.20275e-18
c182 136:14 128:c  c=3.86848e-17
c181 136:14 107:c  c=3.44927e-18
c180 136:14 108:c  c=2.29353e-18
c179 136:14 73:c  c=3.11589e-18
c178 136:14 88:c  c=2.91101e-17
c177 136:14 126:c  c=2.28705e-18
c176 x32|src 61:d  c=5.67946e-19
c175 x32|src 71:d  c=5.67946e-19
c174 x32|src 64:d  c=5.67946e-19
c173 x32|src 56:d  c=2.3592e-18
c172 x32|src 32:rn  c=2.53532e-19
c171 x32|src 53:d  c=5.67946e-19
cg170 135:14 gnd  c=7.3969e-18
c169 135:14 133:c  c=4.07156e-19
c168 135:14 66:d  c=2.36818e-18
c167 135:14 56:d  c=5.49618e-18
c166 135:14 58:d  c=1.65297e-19
c165 135:14 128:c  c=3.31167e-18
c164 135:14 60:d  c=3.004e-18
c163 135:14 54:d  c=2.9639e-19
c162 135:14 130:c  c=3.28693e-18
c161 135:14 109:c  c=2.16454e-18
c160 135:14 116:c  c=2.98128e-18
c159 135:14 88:c  c=2.67776e-18
c158 135:14 65:d  c=3.53734e-18
c157 x26|src 133:c  c=9.73775e-20
c156 x26|src 74:c  c=4.0729e-20
c155 x26|src 82:c  c=1.29384e-20
c154 x26|src 32:rn  c=1.52697e-19
c153 x26|src 60:d  c=5.67946e-19
c152 x26|src 130:c  c=5.57476e-19
c151 x26|src 116:c  c=5.57476e-19
c150 x26|src 126:c  c=1.49779e-20
c149 x26|src 65:d  c=5.67946e-19
c148 x24|drn 82:c  c=7.14964e-21
c147 x24|drn 32:rn  c=1.06443e-20
c146 x24|drn 125:c  c=5.57428e-19
c145 x24|drn 128:c  c=3.17189e-18
c144 x24|drn 107:c  c=5.63452e-19
c143 x24|drn 73:c  c=5.63452e-19
c142 x2|drn 56:d  c=4.3962e-20
c141 x2|drn 57:d  c=5.67946e-19
c140 x2|drn 69:d  c=5.67946e-19
cg139 134:c gnd  c=3.13797e-17
c138 134:c 52:rn  c=8.6749e-17
c137 134:c 32:rn  c=7.86632e-18
cg136 133:c gnd  c=1.25778e-17
c135 133:c 32:rn  c=1.1565e-17
cg134 132:c gnd  c=1.25257e-17
c133 132:c x9|drn  c=1.33078e-19
c132 132:c 50:rn  c=1.40656e-17
cg131 131:c gnd  c=7.02781e-18
c130 131:c 32:rn  c=5.08581e-18
cg129 130:c gnd  c=3.25126e-17
cg128 128:c gnd  c=9.39136e-17
cg127 126:c gnd  c=6.21512e-18
cg126 125:c gnd  c=2.94779e-17
cg125 123:c gnd  c=5.88182e-19
c124 123:c 5:rn  c=2.51143e-20
c123 123:c 41:rn  c=1.0107e-21
c122 122:c 5:rn  c=8.28656e-22
cg121 121:c gnd  c=2.9457e-18
c120 121:c 39:rn  c=3.93379e-21
c119 121:c 5:rn  c=2.2828e-22
c118 121:c 37:rn  c=1.01257e-19
cg117 120:c gnd  c=3.31076e-18
c116 120:c 5:rn  c=1.79183e-20
c115 120:c 41:rn  c=3.50087e-21
cg114 119:c gnd  c=2.28979e-17
cg113 118:c gnd  c=3.05528e-17
c112 118:c 50:rn  c=3.23495e-16
cg111 116:c gnd  c=1.59424e-17
cg110 111:c gnd  c=9.29855e-19
cg109 109:c gnd  c=4.33529e-18
cg108 108:c gnd  c=3.82984e-18
cg107 107:c gnd  c=2.68126e-17
cg106 106:c gnd  c=4.30081e-18
c105 105:c 46:rn  c=1.39252e-17
c104 105:c 43:rn  c=2.87149e-21
cg103 104:c gnd  c=2.94574e-18
c102 104:c 51:rn  c=7.57007e-19
c101 104:c 43:rn  c=1.1823e-19
c100 104:c 41:rn  c=1.43613e-17
cg99 103:c gnd  c=3.91882e-17
c98 103:c 50:rn  c=2.12583e-19
cg97 102:c gnd  c=1.8632e-18
cg96 89:c gnd  c=1.81551e-17
c95 89:c 5:rn  c=3.50496e-19
c94 89:c 41:rn  c=4.38438e-19
cg93 88:c gnd  c=2.6154e-17
c92 88:c 32:rn  c=4.25167e-19
cg91 87:c gnd  c=1.87213e-17
c90 87:c 39:rn  c=1.43055e-17
c89 87:c 37:rn  c=9.76055e-21
cg88 86:c gnd  c=5.67858e-18
c87 86:c 41:rn  c=4.1922e-20
cg86 84:c gnd  c=1.21676e-17
c85 84:c 41:rn  c=3.14415e-20
cg84 83:c gnd  c=1.5947e-17
c83 83:c 52:rn  c=8.09038e-18
c82 83:c 20:rn  c=3.79964e-18
c81 83:c 32:rn  c=8.93125e-17
c80 82:c 1:rn  c=4.88918e-18
c79 82:c 12:rn  c=9.54822e-19
c78 82:c 31:rn  c=5.50732e-18
c77 82:c 51:rn  c=1.36196e-17
c76 82:c x6|src  c=4.86974e-20
c75 82:c 5:rn  c=4.25167e-19
c74 82:c 32:rn  c=1.26788e-15
c73 82:c 41:rn  c=4.25167e-19
c72 82:c 50:rn  c=3.8119e-19
cg71 81:c gnd  c=1.52195e-17
c70 81:c 32:rn  c=8.76674e-17
cg69 77:c gnd  c=2.69804e-17
c68 77:c 39:rn  c=5.80434e-20
c67 77:c 37:rn  c=1.95892e-20
cg66 76:c gnd  c=1.39573e-17
c65 76:c x9|drn  c=3.08189e-20
c64 76:c 50:rn  c=9.58653e-17
cg63 75:c gnd  c=5.76016e-18
c62 75:c x9|drn  c=1.54335e-19
cg61 74:c gnd  c=3.16222e-18
c60 74:c 32:rn  c=9.24426e-17
cg59 73:c gnd  c=1.2181e-17
cg58 72:d gnd  c=3.57636e-17
c57 72:d 52:rn  c=1.0067e-16
c56 72:d 20:rn  c=1.89989e-17
cg55 71:d gnd  c=8.59805e-18
cg54 69:d gnd  c=6.61375e-18
cg53 66:d gnd  c=5.09855e-19
cg52 65:d gnd  c=1.29348e-17
cg51 64:d gnd  c=4.95432e-18
cg50 61:d gnd  c=7.89468e-18
cg49 60:d gnd  c=7.55111e-18
cg48 59:d gnd  c=7.89883e-18
c47 59:d 52:rn  c=5.90592e-18
cg46 58:d gnd  c=1.78258e-17
c45 58:d 52:rn  c=2.87236e-18
cg44 57:d gnd  c=7.33617e-17
c43 57:d 52:rn  c=8.8136e-18
c42 57:d 32:rn  c=2.12583e-19
cg41 56:d gnd  c=2.73286e-17
cg40 54:d gnd  c=3.68675e-18
cg39 53:d gnd  c=3.98892e-18
cg38 52:rn gnd  c=1.49593e-17
cg37 51:rn gnd  c=8.74609e-18
c36 51:rn x6|src  c=7.56515e-20
c35 51:rn m7|x1|drn  c=1.205e-19
cg34 50:rn gnd  c=7.825e-17
c33 50:rn x9|drn  c=1.20946e-19
cg32 49:rn gnd  c=9.42868e-18
cg31 48:rn gnd  c=3.91441e-18
cg30 45:rn gnd  c=6.36768e-18
cg29 44:rn gnd  c=2.87563e-18
cg28 43:rn gnd  c=1.57462e-17
c27 43:rn m7|x1|drn  c=1.50413e-20
cg26 41:rn gnd  c=1.80462e-17
cg25 40:rn gnd  c=6.01717e-18
cg24 39:rn gnd  c=1.92813e-18
cg23 37:rn gnd  c=1.57622e-18
cg22 33:rn gnd  c=8.1721e-18
cg21 32:rn gnd  c=9.53211e-17
c20 32:rn m7|x1|drn  c=4.82645e-20
c19 32:rn x6|src  c=4.79163e-20
cg18 31:rn gnd  c=1.01981e-17
cg17 25:rn gnd  c=4.17871e-18
cg16 23:rn gnd  c=8.1721e-18
cg15 22:rn gnd  c=3.5018e-18
cg14 20:rn gnd  c=1.96921e-17
cg13 12:rn gnd  c=2.02636e-17
cg12 8:rn gnd  c=5.7077e-18
cg11 6:rn gnd  c=7.88627e-18
cg10 5:rn gnd  c=2.15293e-17
cg9 4:rn gnd  c=2.0418e-17
cg8 3:rn gnd  c=3.5018e-18
cg7 2:rn gnd  c=2.57717e-18
cg6 1:rn gnd  c=7.12828e-18
cg5 x9|drn gnd  c=1.01849e-20
cg4 m18|x1|drn gnd  c=6.79162e-20
cg3 x4|src gnd  c=1.23138e-19
cg2 m7|x1|drn gnd  c=1.16777e-19
cg1 x6|src gnd  c=2.89637e-20
r736 530:vdd 531:vdd  r=0.0409063
r735 530:vdd x30|src  r=7.5
r734 527:vdd 529:vdd  r=0.128734
r733 vdd 529:vdd  r=0.109484
r732 vdd 530:vdd  r=0.221375
r731 525:vdd 528:vdd  r=0.0409063
r730 523:vdd 524:vdd  r=0.0409063
r729 523:vdd x29|src  r=7.5
r728 520:vdd 521:vdd  r=0.0409063
r727 518:vdd 522:vdd  r=0.123922
r726 517:vdd 519:vdd  r=0.122719
r725 516:vdd 517:vdd  r=0.181672
r724 514:vdd 515:vdd  r=0.0409063
r723 512:vdd 516:vdd  r=0.129938
r722 511:vdd 513:vdd  r=0.129938
r721 510:vdd 511:vdd  r=0.181672
r720 509:vdd 510:vdd  r=0.123922
r719 508:vdd 509:vdd  r=0.123922
r718 507:vdd 508:vdd  r=0.122719
r717 506:vdd 507:vdd  r=0.122719
r716 505:vdd 506:vdd  r=0.122719
r715 503:vdd x22|src  r=7.5
r714 503:vdd 504:vdd  r=0.0409063
r713 500:vdd 502:vdd  r=0.0409063
r712 498:vdd 499:vdd  r=0.0409063
r711 497:vdd 532:vdd  r=0.0637657
r710 495:vdd 532:vdd  r=0.0601563
r709 494:vdd 501:vdd  r=0.122719
r708 491:vdd 492:vdd  r=0.135953
r707 489:vdd 490:vdd  r=0.0409063
r706 489:vdd x15|src  r=7.5
r705 486:vdd 487:vdd  r=0.0409063
r704 483:vdd 488:vdd  r=0.123922
r703 482:vdd 485:vdd  r=0.0409063
r702 482:vdd 484:vdd  r=0.122719
r701 481:vdd 496:vdd  r=0.0409063
r700 x17|src 481:vdd  r=7.5
r699 480:vdd 484:vdd  r=0.0890313
r698 480:vdd 486:vdd  r=0.221375
r697 480:vdd 483:vdd  r=0.156406
r696 479:vdd 500:vdd  r=0.221375
r695 479:vdd 501:vdd  r=0.17325
r694 478:vdd 493:vdd  r=0.0409063
r693 478:vdd x16|drn  r=7.5
r692 477:vdd 492:vdd  r=0.179266
r691 477:vdd 478:vdd  r=0.206938
r690 476:vdd 526:vdd  r=0.110688
r689 476:vdd 525:vdd  r=0.221375
r688 476:vdd 527:vdd  r=0.146781
r687 475:vdd 503:vdd  r=0.221375
r686 475:vdd 505:vdd  r=0.19611
r685 475:vdd 479:vdd  r=0.385
r684 474:vdd 497:vdd  r=0.156406
r683 474:vdd 498:vdd  r=0.221375
r682 474:vdd 494:vdd  r=0.0890313
r681 473:vdd 491:vdd  r=0.200922
r680 473:vdd 488:vdd  r=0.104672
r679 473:vdd 489:vdd  r=0.221375
r678 472:vdd 519:vdd  r=0.0890313
r677 472:vdd 520:vdd  r=0.221375
r676 472:vdd 518:vdd  r=0.156406
r675 x31|src 525:vdd  r=7.5
r674 x31|src x32|drn  r=0.001
r673 471:vdd 513:vdd  r=0.274313
r672 471:vdd 514:vdd  r=0.206938
r671 471:vdd 512:vdd  r=0.0818126
r670 470:vdd 526:vdd  r=0.878282
r669 470:vdd 522:vdd  r=0.104672
r668 470:vdd 523:vdd  r=0.221375
r667 x27|drn 520:vdd  r=7.5
r666 x27|drn x28|src  r=0.001
r665 x23|src 514:vdd  r=7.5
r664 m10|x1|drn x23|src  r=0.001
r663 x20|src 500:vdd  r=7.5
r662 x21|drn x20|src  r=0.001
r661 x18|drn 498:vdd  r=7.5
r660 x19|drn x18|drn  r=0.001
r659 469:vdd 481:vdd  r=0.221375
r658 469:vdd 495:vdd  r=0.104672
r657 469:vdd 477:vdd  r=0.220172
r656 x13|drn 486:vdd  r=7.5
r655 x13|drn x14|src  r=0.001
r654 x13|bulk 517:vdd  r=7.5
r653 x13|bulk 491:vdd  r=7.5
r652 x13|bulk 526:vdd  r=7.5
r651 x13|bulk 519:vdd  r=7.5
r650 x13|bulk 492:vdd  r=7.5
r649 x13|bulk 482:vdd  r=7.5
r648 x13|bulk 510:vdd  r=7.5
r647 x13|bulk 518:vdd  r=7.5
r646 x13|bulk 527:vdd  r=7.5
r645 x13|bulk 511:vdd  r=7.5
r644 x13|bulk 495:vdd  r=7.5
r643 x13|bulk 469:vdd  r=7.5
r642 x13|bulk 513:vdd  r=7.5
r641 x13|bulk 505:vdd  r=7.5
r640 x13|bulk 473:vdd  r=7.5
r639 x13|bulk 484:vdd  r=7.5
r638 x13|bulk 522:vdd  r=7.5
r637 x13|bulk 497:vdd  r=7.5
r636 x13|bulk 529:vdd  r=7.5
r635 x13|bulk 480:vdd  r=7.5
r634 x13|bulk 506:vdd  r=7.5
r633 x13|bulk 474:vdd  r=7.5
r632 x13|bulk 507:vdd  r=7.5
r631 x13|bulk 508:vdd  r=7.5
r630 x13|bulk 512:vdd  r=7.5
r629 x13|bulk 483:vdd  r=7.5
r628 x13|bulk vdd  r=7.5
r627 x13|bulk 494:vdd  r=7.5
r626 x13|bulk 476:vdd  r=7.5
r625 x13|bulk 470:vdd  r=7.5
r624 x13|bulk 472:vdd  r=7.5
r623 x13|bulk 488:vdd  r=7.5
r622 x13|bulk 516:vdd  r=7.5
r621 x13|bulk 501:vdd  r=7.5
r620 x13|bulk 509:vdd  r=7.5
r619 m11|x1|bulk x33|cathode  r=0.001
r618 m11|x1|bulk x9|bulk  r=0.001
r617 m11|x1|bulk m10|x1|bulk  r=0.001
r616 m11|x1|bulk x10|bulk  r=0.001
r615 m11|x1|bulk x11|bulk  r=0.001
r614 m11|x1|bulk x12|bulk  r=0.001
r613 m11|x1|bulk x13|bulk  r=0.001
r612 m11|x1|bulk x14|bulk  r=0.001
r611 m11|x1|bulk x15|bulk  r=0.001
r610 m11|x1|bulk x16|bulk  r=0.001
r609 m11|x1|bulk x17|bulk  r=0.001
r608 m11|x1|bulk x18|bulk  r=0.001
r607 m11|x1|bulk x19|bulk  r=0.001
r606 m11|x1|bulk x20|bulk  r=0.001
r605 m11|x1|bulk x21|bulk  r=0.001
r604 m11|x1|bulk x22|bulk  r=0.001
r603 m11|x1|bulk x23|bulk  r=0.001
r602 m11|x1|bulk x24|bulk  r=0.001
r601 m11|x1|bulk x25|bulk  r=0.001
r600 m11|x1|bulk x26|bulk  r=0.001
r599 m11|x1|bulk x27|bulk  r=0.001
r598 m11|x1|bulk x28|bulk  r=0.001
r597 m11|x1|bulk x29|bulk  r=0.001
r596 m11|x1|bulk x30|bulk  r=0.001
r595 m11|x1|bulk x31|bulk  r=0.001
r594 x32|bulk m11|x1|bulk  r=0.001
r593 466:gnd 467:gnd  r=0.0409063
r592 466:gnd x8|drn  r=7.5
r591 gnd 466:gnd  r=0.206938
r590 465:gnd gnd  r=0.112204
r589 462:gnd 464:gnd  r=0.0409063
r588 462:gnd m5|x1|src  r=7.5
r587 461:gnd 463:gnd  r=0.1155
r586 459:gnd 460:gnd  r=0.0409063
r585 459:gnd x7|drn  r=7.5
r584 457:gnd 458:gnd  r=0.135953
r583 456:gnd 457:gnd  r=0.359975
r582 455:gnd 456:gnd  r=0.1155
r581 454:gnd 455:gnd  r=0.1155
r580 453:gnd 454:gnd  r=0.571244
r579 452:gnd 453:gnd  r=0.126328
r578 448:gnd 468:gnd  r=0.180469
r577 448:gnd 449:gnd  r=0.135953
r576 445:gnd m23|x1|src  r=7.5
r575 445:gnd 447:gnd  r=0.0409063
r574 443:gnd 446:gnd  r=0.1155
r573 443:gnd 444:gnd  r=0.0409063
r572 442:gnd 450:gnd  r=0.0409063
r571 442:gnd x3|src  r=7.5
r570 441:gnd 468:gnd  r=1.28614
r569 441:gnd 446:gnd  r=0.0962501
r568 441:gnd 445:gnd  r=0.206938
r567 440:gnd 451:gnd  r=0.0433125
r566 440:gnd x4|drn  r=7.5
r565 439:gnd 442:gnd  r=0.206938
r564 439:gnd 449:gnd  r=0.179266
r563 438:gnd 440:gnd  r=0.231
r562 438:gnd 439:gnd  r=0.208141
r561 438:gnd 452:gnd  r=0.169641
r560 437:gnd 465:gnd  r=1.26328
r559 437:gnd 463:gnd  r=0.0962501
r558 437:gnd 462:gnd  r=0.206938
r557 x2|bulk 465:gnd  r=7.5
r556 x2|bulk gnd  r=7.5
r555 m7|x1|bulk 458:gnd  r=7.5
r554 m7|x1|bulk 457:gnd  r=7.5
r553 m5|x1|bulk 463:gnd  r=7.5
r552 m5|x1|bulk 461:gnd  r=7.5
r551 m5|x1|bulk 437:gnd  r=7.5
r550 m23|x1|bulk 446:gnd  r=7.5
r549 m23|x1|bulk 443:gnd  r=7.5
r548 m23|x1|bulk 441:gnd  r=7.5
r547 m18|x1|bulk x4|bulk  r=0.001
r546 m18|x1|bulk x5|bulk  r=0.001
r545 m18|x1|bulk x6|bulk  r=0.001
r544 m18|x1|bulk x7|bulk  r=0.001
r543 m18|x1|bulk x8|bulk  r=0.001
r542 m18|x1|bulk m23|x1|bulk  r=0.001
r541 m18|x1|bulk m5|x1|bulk  r=0.001
r540 m18|x1|bulk 448:gnd  r=7.5
r539 m18|x1|bulk m7|x1|bulk  r=0.001
r538 m18|x1|bulk x1|bulk  r=0.001
r537 m18|x1|bulk 449:gnd  r=7.5
r536 m18|x1|bulk 452:gnd  r=7.5
r535 m18|x1|bulk 453:gnd  r=7.5
r534 m18|x1|bulk x2|bulk  r=0.001
r533 m18|x1|bulk x3|bulk  r=0.001
r532 x33|anode 456:gnd  r=7.5
r531 x33|anode 455:gnd  r=7.5
r530 x33|anode 454:gnd  r=7.5
r529 x33|anode m18|x1|bulk  r=0.001
r528 436:gnd 461:gnd  r=0.585922
r527 436:gnd 458:gnd  r=0.282735
r526 436:gnd 459:gnd  r=0.206938
r525 433:3 m10|x1|src  r=7.5
r524 433:3 3  r=0.03675
r523 431:3 432:3  r=0.037625
r522 429:3 434:3  r=0.04025
r521 429:3 431:3  r=0.002625
r520 428:3 430:3  r=0.0405238
r519 428:3 429:3  r=4.5
r518 426:3 427:3  r=0.282434
r517 426:3 428:3  r=0.0405238
r516 424:3 427:3  r=0.0405238
r515 424:3 425:3  r=0.0405238
r514 423:3 435:3  r=0.04025
r513 423:3 433:3  r=0.0035
r512 423:3 424:3  r=4.5
r511 m11|x1|drn 431:3  r=7.5
r510 x23|drn m11|x1|drn  r=0.001
r509 412:cn 413:cn  r=11.4286
r508 409:cn 410:cn  r=7.85716
r507 407:cn 408:cn  r=1.57558
r506 403:cn 416:cn  r=27.6786
r505 402:cn 404:cn  r=2.64833
r504 402:cn 403:cn  r=2.64707
r503 401:cn 421:cn  r=0.039375
r502 401:cn 402:cn  r=7.5
r501 399:cn 420:cn  r=0.039375
r500 397:cn 418:cn  r=0.039375
r499 395:cn 419:cn  r=0.039375
r498 x2|gate 416:cn  r=3.92858
r497 394:cn 417:cn  r=7.85716
r496 394:cn x2|gate  r=3.92858
r495 x12|gate 393:cn  r=3.92858
r494 392:cn 415:cn  r=11.4286
r493 392:cn x12|gate  r=3.92858
r492 x11|gate 391:cn  r=3.92858
r491 390:cn x11|gate  r=3.92858
r490 390:cn 414:cn  r=11.4286
r489 x10|gate 412:cn  r=3.92858
r488 389:cn x10|gate  r=3.92858
r487 m18|x1|gate 410:cn  r=3.92858
r486 388:cn 411:cn  r=7.85716
r485 388:cn m18|x1|gate  r=3.92858
r484 386:cn 405:cn  r=2.95692
r483 384:cn 401:cn  r=0.000875001
r482 384:cn 385:cn  r=0.04025
r481 383:cn 386:cn  r=0.0405238
r480 383:cn 384:cn  r=4.5
r479 380:cn 399:cn  r=0.000875001
r478 380:cn 381:cn  r=0.04025
r477 379:cn 405:cn  r=0.0374066
r476 379:cn 382:cn  r=0.0374066
r475 379:cn 380:cn  r=4.5
r474 376:cn 397:cn  r=0.000875001
r473 376:cn 377:cn  r=0.04025
r472 375:cn 378:cn  r=0.0405238
r471 375:cn 376:cn  r=4.5
r470 373:cn 395:cn  r=0.000875001
r469 373:cn 374:cn  r=0.04025
r468 372:cn 407:cn  r=0.0528572
r467 372:cn 373:cn  r=4.5
r466 371:cn 400:cn  r=3.50001
r465 371:cn 399:cn  r=7.5
r464 370:cn 371:cn  r=2.00001
r463 369:cn 398:cn  r=3.50001
r462 369:cn 397:cn  r=7.5
r461 368:cn 369:cn  r=3.50001
r460 367:cn 389:cn  r=10.3572
r459 367:cn 368:cn  r=79.4645
r458 366:cn 396:cn  r=3.50001
r457 366:cn 395:cn  r=7.5
r456 365:cn 366:cn  r=2.58774
r455 365:cn 409:cn  r=21.7858
r454 363:cn 383:cn  r=0.0405238
r453 363:cn 364:cn  r=0.530334
r452 362:cn 378:cn  r=1.19788
r451 362:cn 372:cn  r=0.0405238
r450 360:cn 406:cn  r=7.85716
r449 m11|x1|gate 361:cn  r=3.92858
r448 m11|x1|gate 360:cn  r=3.92858
r447 359:cn 367:cn  r=21.9347
r446 359:cn 391:cn  r=10.3572
r445 358:cn 387:cn  r=0.0405238
r444 358:cn 364:cn  r=0.0405238
r443 357:cn 422:cn  r=0.04025
r442 357:cn cn  r=0.0279125
r441 357:cn 358:cn  r=4.5
r440 356:cn 359:cn  r=21.9347
r439 356:cn 393:cn  r=10.3572
r438 355:cn 382:cn  r=0.729209
r437 355:cn 375:cn  r=0.0405238
r436 354:cn 361:cn  r=101.25
r435 354:cn 370:cn  r=13.2143
r434 345:2 346:2  r=0.357144
r433 m5|x1|gate 346:2  r=3.92858
r432 342:2 m5|x1|gate  r=3.92858
r431 342:2 2  r=7.85716
r430 341:2 345:2  r=69.643
r429 340:2 344:2  r=11.4286
r428 339:2 343:2  r=11.4286
r427 x27|gate 339:2  r=3.92858
r426 336:2 x27|gate  r=3.92858
r425 335:2 353:2  r=0.039375
r424 333:2 337:2  r=0.0402907
r423 333:2 334:2  r=0.0402907
r422 331:2 332:2  r=0.0409063
r421 331:2 348:2  r=0.770001
r420 329:2 330:2  r=0.035
r419 x29|gate 328:2  r=3.92858
r418 327:2 351:2  r=11.4286
r417 327:2 x29|gate  r=3.92858
r416 x28|gate 340:2  r=3.92858
r415 326:2 x28|gate  r=3.92858
r414 325:2 336:2  r=11.4286
r413 322:2 338:2  r=0.17325
r412 322:2 323:2  r=0.0409063
r411 321:2 349:2  r=0.724282
r410 321:2 324:2  r=0.0409063
r409 318:2 352:2  r=0.04025
r408 318:2 329:2  r=0.00525001
r407 317:2 320:2  r=0.0405238
r406 317:2 319:2  r=0.0405238
r405 317:2 318:2  r=4.5
r404 315:2 350:2  r=0.0405238
r403 312:2 315:2  r=4.5
r402 312:2 347:2  r=0.04025
r401 312:2 316:2  r=0.04025
r400 311:2 337:2  r=0.205735
r399 311:2 348:2  r=0.535391
r398 311:2 347:2  r=0.366953
r397 310:2 338:2  r=0.0542501
r396 310:2 349:2  r=0.163625
r395 309:2 341:2  r=2.81251
r394 309:2 333:2  r=7.5
r393 308:2 309:2  r=2.81251
r392 x24|src 312:2  r=7.5
r391 307:2 320:2  r=0.283667
r390 307:2 315:2  r=0.0405238
r389 304:2 305:2  r=1.68243
r388 304:2 310:2  r=4.5
r387 304:2 313:2  r=0.0551298
r386 x2|src 331:2  r=7.5
r385 303:2 328:2  r=11.4286
r384 301:2 335:2  r=7.5
r383 301:2 302:2  r=3.50001
r382 300:2 301:2  r=3.50001
r381 m7|x1|src 321:2  r=7.5
r380 299:2 306:2  r=0.037
r379 299:2 305:2  r=0.037
r378 298:2 335:2  r=0.000875001
r377 298:2 314:2  r=0.04025
r376 298:2 299:2  r=4.5
r375 297:2 303:2  r=16.6072
r374 297:2 308:2  r=21.2501
r373 297:2 300:2  r=12.8572
r372 296:2 326:2  r=11.4286
r371 296:2 303:2  r=28.5715
r370 296:2 325:2  r=28.5715
r369 x25|drn 329:2  r=7.5
r368 x26|drn x25|drn  r=0.001
r367 m11|x1|src 322:2  r=7.5
r366 286:4 288:4  r=68.2145
r365 285:4 290:4  r=0.635251
r364 x4|gate 288:4  r=7.85716
r363 284:4 x4|gate  r=7.85716
r362 284:4 4  r=7.85716
r361 283:4 287:4  r=15.3572
r360 278:4 280:4  r=11.4286
r359 275:4 287:4  r=3.15001
r358 275:4 286:4  r=3.15001
r357 274:4 295:4  r=0.0402907
r356 274:4 275:4  r=7.5
r355 272:4 290:4  r=0.0402907
r354 272:4 273:4  r=0.0402907
r353 270:4 291:4  r=0.0507577
r352 269:4 271:4  r=0.039375
r351 x19|gate 276:4  r=3.92858
r350 268:4 292:4  r=11.4286
r349 268:4 x19|gate  r=3.92858
r348 x18|gate 267:4  r=3.92858
r347 266:4 282:4  r=11.4286
r346 266:4 x18|gate  r=3.92858
r345 264:4 265:4  r=0.0409063
r344 x17|gate 278:4  r=3.92858
r343 263:4 281:4  r=10.3572
r342 263:4 x17|gate  r=3.92858
r341 261:4 262:4  r=0.0409063
r340 258:4 293:4  r=0.04025
r339 258:4 269:4  r=0.000875001
r338 257:4 260:4  r=0.0405239
r337 257:4 259:4  r=0.0405239
r336 257:4 258:4  r=4.5
r335 256:4 294:4  r=0.0405239
r334 253:4 277:4  r=0.0405238
r333 253:4 254:4  r=0.0405238
r332 252:4 289:4  r=0.04025
r331 252:4 256:4  r=4.5
r330 252:4 255:4  r=0.04025
r329 251:4 291:4  r=0.559237
r328 250:4 274:4  r=0.0273082
r327 249:4 261:4  r=0.972126
r326 x10|src 252:4  r=7.5
r325 x9|src 261:4  r=7.5
r324 248:4 279:4  r=3.50001
r323 248:4 272:4  r=7.5
r322 247:4 248:4  r=3.50001
r321 246:4 260:4  r=0.2849
r320 246:4 256:4  r=0.0405239
r319 m18|x1|src 264:4  r=7.5
r318 x1|drn 270:4  r=7.5
r317 245:4 281:4  r=21.9347
r316 245:4 267:4  r=10.3572
r315 244:4 276:4  r=10.3572
r314 244:4 245:4  r=21.8626
r313 243:4 244:4  r=16.0715
r312 243:4 247:4  r=71.4287
r311 243:4 283:4  r=70.5359
r310 x11|drn 269:4  r=7.5
r309 x12|drn x11|drn  r=0.001
r308 242:4 289:4  r=0.300782
r307 242:4 250:4  r=0.416291
r306 242:4 251:4  r=0.386814
r305 241:4 253:4  r=4.5
r304 241:4 249:4  r=0.449969
r303 241:4 264:4  r=0.401844
r302 241:4 285:4  r=0.0560001
r301 233:9 234:9  r=16.7858
r300 231:9 9  r=7.85716
r299 230:9 232:9  r=22.8572
r298 227:9 234:9  r=3.50001
r297 227:9 228:9  r=3.50001
r296 226:9 238:9  r=0.039375
r295 226:9 227:9  r=7.5
r294 224:9 232:9  r=3.38711
r293 224:9 225:9  r=3.38711
r292 223:9 237:9  r=0.0402907
r291 223:9 224:9  r=7.5
r290 221:9 222:9  r=0.0409063
r289 220:9 240:9  r=0.0409063
r288 218:9 219:9  r=0.0409063
r287 216:9 x12|src  r=7.5
r286 216:9 239:9  r=0.0409063
r285 215:9 217:9  r=0.04025
r284 215:9 x1|src  r=7.5
r283 215:9 235:9  r=0.04025
r282 210:9 226:9  r=0.000875001
r281 210:9 211:9  r=0.04025
r280 209:9 213:9  r=0.0405238
r279 209:9 212:9  r=0.0405238
r278 209:9 210:9  r=4.5
r277 x7|gate 231:9  r=3.92858
r276 208:9 214:9  r=0.0409063
r275 207:9 220:9  r=0.216563
r274 207:9 221:9  r=0.741126
r273 206:9 223:9  r=0.0402907
r272 205:9 216:9  r=0.216563
r271 205:9 235:9  r=0.685782
r270 204:9 x7|gate  r=3.92858
r269 203:9 204:9  r=19.4643
r268 203:9 233:9  r=50.0001
r267 203:9 225:9  r=79.1073
r266 202:9 205:9  r=0.385
r265 202:9 208:9  r=0.216563
r264 201:9 236:9  r=0.0405238
r263 201:9 215:9  r=4.5
r262 200:9 201:9  r=0.0405238
r261 200:9 213:9  r=0.958548
r260 x27|src 218:9  r=7.5
r259 199:9 229:9  r=7.85716
r258 m10|x1|gate 230:9  r=3.92858
r257 m10|x1|gate 199:9  r=3.92858
r256 x28|drn 220:9  r=7.5
r255 x29|drn x28|drn  r=0.001
r254 198:9 218:9  r=0.216563
r253 198:9 206:9  r=0.229797
r252 198:9 207:9  r=0.385
r251 x10|drn 208:9  r=7.5
r250 x11|src x10|drn  r=0.001
r249 m5|x1|drn 221:9  r=7.5
r248 196:q 197:q  r=0.0409063
r247 193:q 195:q  r=0.0409063
r246 192:q 194:q  r=0.0409063
r245 191:q 193:q  r=0.463204
r244 191:q q  r=0.170122
r243 m23|x1|drn 193:q  r=7.5
r242 x13|src 192:q  r=7.5
r241 190:q 196:q  r=0.218969
r240 x14|drn x15|drn  r=0.001
r239 x14|drn 196:q  r=7.5
r238 189:q 190:q  r=0.385
r237 189:q 192:q  r=0.218969
r236 189:q 191:q  r=0.275516
r235 186:16 187:16  r=0.567876
r234 185:16 16  r=7.85716
r233 x16|gate 182:16  r=3.92858
r232 181:16 188:16  r=7.85716
r231 181:16 x16|gate  r=3.92858
r230 176:16 186:16  r=0.282735
r229 175:16 184:16  r=2.31334
r228 175:16 183:16  r=3.50001
r227 174:16 176:16  r=0.0402907
r226 174:16 175:16  r=7.5
r225 171:16 172:16  r=0.0409063
r224 169:16 170:16  r=0.0409063
r223 167:16 168:16  r=0.0409063
r222 x15|gate 166:16  r=3.92858
r221 165:16 180:16  r=11.4286
r220 165:16 x15|gate  r=3.92858
r219 x14|gate 164:16  r=3.92858
r218 163:16 179:16  r=11.4286
r217 163:16 x14|gate  r=3.92858
r216 162:16 178:16  r=7.85716
r215 m23|x1|gate 162:16  r=3.92858
r214 161:16 m23|x1|gate  r=3.92858
r213 x13|gate 160:16  r=3.92858
r212 159:16 177:16  r=11.4286
r211 159:16 x13|gate  r=3.92858
r210 158:16 x5|drn  r=7.5
r209 158:16 187:16  r=0.222578
r208 158:16 173:16  r=0.0433125
r207 157:16 167:16  r=0.216563
r206 156:16 174:16  r=0.0402907
r205 x3|gate 185:16  r=3.92858
r204 155:16 183:16  r=75.1788
r203 155:16 x3|gate  r=3.92858
r202 154:16 161:16  r=6.07144
r201 153:16 154:16  r=29.1072
r200 152:16 160:16  r=10.3572
r199 152:16 153:16  r=86.9645
r198 151:16 171:16  r=0.216563
r197 150:16 153:16  r=150.893
r196 149:16 150:16  r=55.0001
r195 149:16 184:16  r=110
r194 148:16 152:16  r=21.9347
r193 148:16 164:16  r=10.3572
r192 147:16 151:16  r=0.385
r191 147:16 157:16  r=0.354321
r190 147:16 169:16  r=0.216563
r189 147:16 156:16  r=0.103469
r188 146:16 182:16  r=46.2501
r187 146:16 149:16  r=17.1429
r186 x21|src 171:16  r=7.5
r185 x22|drn x21|src  r=0.001
r184 x19|src 169:16  r=7.5
r183 x20|drn x19|src  r=0.001
r182 x17|drn 167:16  r=7.5
r181 x17|drn x18|src  r=0.001
r180 145:16 148:16  r=21.9347
r179 145:16 166:16  r=10.3572
r178 143:14 144:14  r=0.0409063
r177 142:14 14  r=0.0409063
r176 140:14 141:14  r=0.0409063
r175 138:14 139:14  r=0.0409063
r174 137:14 143:14  r=0.218969
r173 137:14 142:14  r=0.738719
r172 136:14 138:14  r=0.218969
r171 x32|src 143:14  r=7.5
r170 x32|src x30|drn  r=0.001
r169 135:14 140:14  r=0.218969
r168 135:14 137:14  r=0.385
r167 135:14 136:14  r=0.385
r166 x26|src 140:14  r=7.5
r165 x26|src x31|drn  r=0.001
r164 x24|drn 138:14  r=7.5
r163 x25|src x24|drn  r=0.001
r162 x2|drn 142:14  r=7.5
r161 x8|src x2|drn  r=0.001
r160 125:c 127:c  r=11.4286
r159 x1|gate 122:c  r=3.92858
r158 121:c x1|gate  r=3.92858
r157 120:c 122:c  r=6.60716
r156 120:c 123:c  r=1.24408
r155 114:c 126:c  r=3.50001
r154 114:c 115:c  r=3.50001
r153 113:c 133:c  r=0.039375
r152 113:c 114:c  r=7.5
r151 112:c 131:c  r=0.039375
r150 110:c 132:c  r=0.039375
r149 x26|gate 116:c  r=3.92858
r148 109:c 130:c  r=11.4286
r147 109:c x26|gate  r=3.92858
r146 x25|gate 108:c  r=3.92858
r145 107:c x25|gate  r=3.92858
r144 107:c 129:c  r=11.4286
r143 x24|gate 125:c  r=3.92858
r142 106:c 128:c  r=11.4286
r141 106:c x24|gate  r=3.92858
r140 m7|x1|gate 105:c  r=3.92858
r139 104:c 124:c  r=7.85716
r138 104:c m7|x1|gate  r=3.92858
r137 x9|gate 103:c  r=3.92858
r136 102:c 119:c  r=7.85716
r135 102:c x9|gate  r=3.92858
r134 99:c 113:c  r=0.000875001
r133 99:c 100:c  r=0.04025
r132 98:c 101:c  r=0.0405238
r131 98:c 99:c  r=4.5
r130 97:c 118:c  r=2.21229
r129 95:c 112:c  r=0.000875001
r128 95:c 96:c  r=0.04025
r127 94:c 97:c  r=0.0405238
r126 94:c 95:c  r=4.5
r125 93:c 117:c  r=0.592001
r124 91:c 110:c  r=0.000875001
r123 91:c 92:c  r=0.04025
r122 90:c 93:c  r=0.0405239
r121 90:c 91:c  r=4.5
r120 89:c 123:c  r=51.0716
r119 88:c 116:c  r=11.4286
r118 88:c 126:c  r=56.4287
r117 87:c 105:c  r=10.3572
r116 85:c 112:c  r=7.5
r115 85:c 86:c  r=3.50001
r114 84:c 89:c  r=31.2501
r113 84:c 85:c  r=3.50001
r112 81:c 94:c  r=0.0405238
r111 81:c 101:c  r=2.55917
r110 80:c 111:c  r=3.50001
r109 80:c 110:c  r=7.5
r108 79:c 83:c  r=0.0405238
r107 79:c 82:c  r=0.0405238
r106 78:c 134:c  r=0.04025
r105 78:c c  r=0.02135
r104 78:c 79:c  r=4.5
r103 77:c 121:c  r=10.3572
r102 77:c 87:c  r=87.079
r101 76:c 90:c  r=0.0405239
r100 76:c 118:c  r=0.803209
r99 75:c 80:c  r=4.54374
r98 75:c 103:c  r=72.5002
r97 74:c 98:c  r=0.0405238
r96 74:c 82:c  r=0.969709
r95 73:c 128:c  r=28.5715
r94 73:c 108:c  r=11.4286
r93 73:c 88:c  r=28.5715
r92 69:d 70:d  r=7.85716
r91 x31|gate 66:d  r=3.92858
r90 65:d 67:d  r=11.4286
r89 65:d x31|gate  r=3.92858
r88 x30|gate 64:d  r=3.92858
r87 63:d 71:d  r=11.4286
r86 63:d x30|gate  r=3.92858
r85 x32|gate 62:d  r=3.92858
r84 61:d 68:d  r=11.4286
r83 61:d x32|gate  r=3.92858
r82 60:d 66:d  r=11.0715
r81 x8|gate 69:d  r=3.92858
r80 57:d x8|gate  r=3.92858
r79 56:d 64:d  r=11.0715
r78 55:d 59:d  r=3.50001
r77 55:d 58:d  r=3.50001
r76 d 72:d  r=0.0603466
r75 d 55:d  r=7.5
r74 54:d 58:d  r=32.1429
r73 54:d 57:d  r=111.072
r72 54:d 56:d  r=12.1429
r71 53:d 62:d  r=11.0715
r70 53:d 56:d  r=28.5715
r69 53:d 60:d  r=28.5715
r68 44:rn 45:rn  r=17.6786
r67 43:rn 44:rn  r=13.2143
r66 41:rn 46:rn  r=78.9288
r65 40:rn 42:rn  r=7.85716
r64 x6|gate 46:rn  r=3.92858
r63 39:rn x6|gate  r=3.92858
r62 39:rn 47:rn  r=7.85716
r61 37:rn 38:rn  r=7.85716
r60 x20|gate 34:rn  r=3.92858
r59 33:rn 35:rn  r=11.4286
r58 33:rn x20|gate  r=3.92858
r57 32:rn 50:rn  r=1.54321
r56 30:rn 45:rn  r=3.50001
r55 30:rn 41:rn  r=3.50001
r54 29:rn 51:rn  r=0.039375
r53 29:rn 30:rn  r=7.5
r52 28:rn 48:rn  r=0.039375
r51 x23|gate 40:rn  r=3.92858
r50 27:rn 43:rn  r=24.8215
r49 27:rn x23|gate  r=3.92858
r48 26:rn 49:rn  r=11.4286
r47 x22|gate 26:rn  r=3.92858
r46 25:rn x22|gate  r=3.92858
r45 x21|gate 24:rn  r=3.92858
r44 23:rn x21|gate  r=3.92858
r43 23:rn 36:rn  r=11.4286
r42 22:rn 34:rn  r=10.3572
r41 21:rn 31:rn  r=3.15425
r40 19:rn 52:rn  r=0.04025
r39 19:rn rn  r=0.0279125
r38 18:rn 21:rn  r=0.0405238
r37 18:rn 20:rn  r=0.0405238
r36 18:rn 19:rn  r=4.5
r35 15:rn 29:rn  r=0.000875001
r34 15:rn 16:rn  r=0.04025
r33 14:rn 31:rn  r=0.0395814
r32 14:rn 17:rn  r=0.0395814
r31 14:rn 15:rn  r=4.5
r30 10:rn 28:rn  r=0.000875001
r29 10:rn 11:rn  r=0.04025
r28 9:rn 13:rn  r=0.0405238
r27 9:rn 12:rn  r=0.0405238
r26 9:rn 10:rn  r=4.5
r25 7:rn 28:rn  r=7.5
r24 7:rn 8:rn  r=3.50001
r23 6:rn 7:rn  r=3.50001
r22 x5|gate 37:rn  r=7.85716
r21 5:rn x5|gate  r=7.85716
r20 4:rn 25:rn  r=10.3572
r19 3:rn 4:rn  r=22.5058
r18 3:rn 22:rn  r=21.9347
r17 3:rn 24:rn  r=10.3572
r16 2:rn 4:rn  r=14.6429
r15 2:rn 5:rn  r=100
r14 2:rn 6:rn  r=12.6786
r13 1:rn 17:rn  r=1.62183
r12 1:rn 32:rn  r=1.10692
r11 1:rn 12:rn  r=0.146458
r10 22 x9|drn  r=0.001
r9 22 x16|src  r=0.001
r8 18 m18|x1|drn  r=0.001
r7 18 x3|drn  r=0.001
r6 20 x4|src  r=0.001
r5 20 x5|src  r=0.001
r4 19 m7|x1|drn  r=0.001
r3 19 x6|drn  r=0.001
r2 21 x6|src  r=0.001
r1 21 x7|src  r=0.001
x9 x9|drn x9|gate x9|src x9|bulk PE w=0.22u l=0.18u as=0.0275p ad=0.1984p ps=0.47u
+  pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x32 x32|drn x32|gate x32|src x32|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x31 x31|drn x31|gate x31|src x31|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x30 x30|drn x30|gate x30|src x30|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1984p
+ ps=1.04u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x29 x29|drn x29|gate x29|src x29|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1984p
+ ps=1.04u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x28 x28|drn x28|gate x28|src x28|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x27 x27|drn x27|gate x27|src x27|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1984p
+ ps=1.04u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x26 x26|drn x26|gate x26|src x26|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x25 x25|drn x25|gate x25|src x25|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x24 x24|drn x24|gate x24|src x24|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1984p
+ ps=1.04u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x23 x23|drn x23|gate x23|src x23|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x22 x22|drn x22|gate x22|src x22|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1984p
+ ps=1.04u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x21 x21|drn x21|gate x21|src x21|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x20 x20|drn x20|gate x20|src x20|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x19 x19|drn x19|gate x19|src x19|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x18 x18|drn x18|gate x18|src x18|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x17 x17|drn x17|gate x17|src x17|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1984p
+ ps=1.04u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x16 x16|drn x16|gate x16|src x16|bulk PE w=0.22u l=0.18u as=0.1984p ad=0.0275p
+ ps=1.88u pd=0.47u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x15 x15|drn x15|gate x15|src x15|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1984p
+ ps=1.04u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x14 x14|drn x14|gate x14|src x14|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x13 x13|drn x13|gate x13|src x13|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1984p
+ ps=1.04u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x12 x12|drn x12|gate x12|src x12|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1984p
+ ps=1.04u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x11 x11|drn x11|gate x11|src x11|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1102p
+ ps=1.04u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x10 x10|drn x10|gate x10|src x10|bulk PE w=0.22u l=0.18u as=0.1102p ad=0.1984p
+ ps=1.04u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
xm11|x1 m11|x1|drn m11|x1|gate m11|x1|src m11|x1|bulk PE w=0.22u l=0.18u as=0.1984p
+  ad=0.1102p ps=1.88u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
xm10|x1 m10|x1|drn m10|x1|gate m10|x1|src m10|x1|bulk PE w=0.22u l=0.18u as=0.1984p
+  ad=0.1102p ps=1.88u pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)'
x8 x8|drn x8|gate x8|src x8|bulk NE w=0.22u l=0.18u as=0.1984p ad=0.1102p ps=1.88u
+  pd=1.04u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
x7 x7|drn x7|gate x7|src x7|bulk NE w=0.22u l=0.18u as=0.1984p ad=0.0275p ps=1.88u
+  pd=0.47u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
x6 x6|drn x6|gate x6|src x6|bulk NE w=0.22u l=0.18u as=0.0275p ad=0.0275p ps=0.47u
+  pd=0.47u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
x5 x5|drn x5|gate x5|src x5|bulk NE w=0.44u l=0.18u as=0.2112p ad=0.055p ps=1.84u
+  pd=0.69u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
x4 x4|drn x4|gate x4|src x4|bulk NE w=0.44u l=0.18u as=0.2112p ad=0.055p ps=1.84u
+  pd=0.69u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
x3 x3|drn x3|gate x3|src x3|bulk NE w=0.22u l=0.18u as=0.1984p ad=0.0275p ps=1.88u
+  pd=0.47u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
x2 x2|drn x2|gate x2|src x2|bulk NE w=0.22u l=0.18u as=0.1102p ad=0.1984p ps=1.04u
+  pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
x1 x1|drn x1|gate x1|src x1|bulk NE w=0.22u l=0.18u as=0.1984p ad=0.1984p ps=1.88u
+  pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
xm7|x1 m7|x1|drn m7|x1|gate m7|x1|src m7|x1|bulk NE w=0.22u l=0.18u as=0.1984p
+ ad=0.0275p ps=1.88u pd=0.47u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
xm5|x1 m5|x1|drn m5|x1|gate m5|x1|src m5|x1|bulk NE w=0.22u l=0.18u as=0.1984p
+ ad=0.1984p ps=1.88u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
xm23|x1 m23|x1|drn m23|x1|gate m23|x1|src m23|x1|bulk NE w=0.22u l=0.18u as=0.1984p
+  ad=0.1984p ps=1.88u pd=1.88u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
xm18|x1 m18|x1|drn m18|x1|gate m18|x1|src m18|x1|bulk NE w=0.22u l=0.18u as=0.1984p
+  ad=0.0275p ps=1.88u pd=0.47u nrs=-1 nrd=-1 m='(1*1)' par1='(1*1)' xf_subext=0
x33 x33|anode x33|cathode dnw area=51.0769p perimeter=58.37u dbv=0.0 m=1
+ xf_subext=0

.ends

